module MuxLookup_Test( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input  [1:0]  io_PC_Sel, // @[:@6.4]
  input  [31:0] io_pc_out, // @[:@6.4]
  input  [31:0] io_pc_recover, // @[:@6.4]
  input  [31:0] io_new_addr, // @[:@6.4]
  output [31:0] io_next_pc, // @[:@6.4]
  output [31:0] io_pc_4 // @[:@6.4]
);
  wire [32:0] _T_18; // @[MuxLookup_Test.scala 18:24:@8.4]
  wire  _T_24; // @[Mux.scala 46:19:@11.4]
  wire [31:0] _T_25; // @[Mux.scala 46:16:@12.4]
  wire  _T_26; // @[Mux.scala 46:19:@13.4]
  wire [31:0] _T_27; // @[Mux.scala 46:16:@14.4]
  wire  _T_28; // @[Mux.scala 46:19:@15.4]
  assign _T_18 = io_pc_out + 32'h4; // @[MuxLookup_Test.scala 18:24:@8.4]
  assign _T_24 = 2'h2 == io_PC_Sel; // @[Mux.scala 46:19:@11.4]
  assign _T_25 = _T_24 ? io_new_addr : 32'h0; // @[Mux.scala 46:16:@12.4]
  assign _T_26 = 2'h1 == io_PC_Sel; // @[Mux.scala 46:19:@13.4]
  assign _T_27 = _T_26 ? io_pc_recover : _T_25; // @[Mux.scala 46:16:@14.4]
  assign _T_28 = 2'h0 == io_PC_Sel; // @[Mux.scala 46:19:@15.4]
  assign io_next_pc = _T_28 ? io_pc_4 : _T_27; // @[MuxLookup_Test.scala 20:14:@17.4]
  assign io_pc_4 = io_pc_out + 32'h4; // @[MuxLookup_Test.scala 18:11:@10.4]
endmodule
