module ALU(
  input         clock,
  input         reset,
  input  [31:0] io_Src_A,
  input  [31:0] io_Src_B,
  input  [4:0]  io_ALUOp,
  output [31:0] io_Sum,
  output        io_Conflag
);
  wire [5:0] shamt; // @[ALU.scala 54:23]
  wire [32:0] _T_32; // @[ALU.scala 56:28]
  wire [31:0] _T_33; // @[ALU.scala 56:28]
  wire [32:0] _T_34; // @[ALU.scala 57:28]
  wire [32:0] _T_35; // @[ALU.scala 57:28]
  wire [31:0] _T_36; // @[ALU.scala 57:28]
  wire [31:0] _T_37; // @[ALU.scala 58:28]
  wire [31:0] _T_38; // @[ALU.scala 59:28]
  wire [31:0] _GEN_0; // @[ALU.scala 60:28]
  wire [31:0] _T_39; // @[ALU.scala 60:28]
  wire [94:0] _GEN_1; // @[ALU.scala 61:28]
  wire [94:0] _T_40; // @[ALU.scala 61:28]
  wire [31:0] _T_41; // @[ALU.scala 62:28]
  wire [31:0] _T_42; // @[ALU.scala 63:34]
  wire [31:0] _T_43; // @[ALU.scala 63:37]
  wire [31:0] _T_44; // @[ALU.scala 63:53]
  wire [31:0] _T_46; // @[ALU.scala 64:54]
  wire  _T_47; // @[ALU.scala 64:37]
  wire  _T_48; // @[ALU.scala 65:28]
  wire  _T_49; // @[Mux.scala 46:19]
  wire [31:0] _T_50; // @[Mux.scala 46:16]
  wire  _T_51; // @[Mux.scala 46:19]
  wire [31:0] _T_52; // @[Mux.scala 46:16]
  wire  _T_53; // @[Mux.scala 46:19]
  wire [31:0] _T_54; // @[Mux.scala 46:16]
  wire  _T_55; // @[Mux.scala 46:19]
  wire [31:0] _T_56; // @[Mux.scala 46:16]
  wire  _T_57; // @[Mux.scala 46:19]
  wire [94:0] _T_58; // @[Mux.scala 46:16]
  wire  _T_59; // @[Mux.scala 46:19]
  wire [94:0] _T_60; // @[Mux.scala 46:16]
  wire  _T_61; // @[Mux.scala 46:19]
  wire [94:0] _T_62; // @[Mux.scala 46:16]
  wire  _T_63; // @[Mux.scala 46:19]
  wire [94:0] _T_64; // @[Mux.scala 46:16]
  wire  _T_65; // @[Mux.scala 46:19]
  wire [94:0] _T_66; // @[Mux.scala 46:16]
  wire  _T_67; // @[Mux.scala 46:19]
  wire [94:0] _T_68; // @[Mux.scala 46:16]
  wire  _T_72; // @[ALU.scala 69:37]
  wire  _T_75; // @[ALU.scala 70:37]
  wire  _T_81; // @[ALU.scala 72:37]
  wire  _T_83; // @[ALU.scala 74:28]
  wire  _T_84; // @[Mux.scala 46:19]
  wire  _T_85; // @[Mux.scala 46:16]
  wire  _T_86; // @[Mux.scala 46:19]
  wire  _T_87; // @[Mux.scala 46:16]
  wire  _T_88; // @[Mux.scala 46:19]
  wire  _T_89; // @[Mux.scala 46:16]
  wire  _T_90; // @[Mux.scala 46:19]
  wire  _T_91; // @[Mux.scala 46:16]
  wire  _T_92; // @[Mux.scala 46:19]
  wire  _T_93; // @[Mux.scala 46:16]
  wire  _T_94; // @[Mux.scala 46:19]
  assign shamt = io_Src_B[5:0]; // @[ALU.scala 54:23]
  assign _T_32 = io_Src_A + io_Src_B; // @[ALU.scala 56:28]
  assign _T_33 = io_Src_A + io_Src_B; // @[ALU.scala 56:28]
  assign _T_34 = io_Src_A - io_Src_B; // @[ALU.scala 57:28]
  assign _T_35 = $unsigned(_T_34); // @[ALU.scala 57:28]
  assign _T_36 = _T_35[31:0]; // @[ALU.scala 57:28]
  assign _T_37 = io_Src_A & io_Src_B; // @[ALU.scala 58:28]
  assign _T_38 = io_Src_A | io_Src_B; // @[ALU.scala 59:28]
  assign _GEN_0 = {{26'd0}, shamt}; // @[ALU.scala 60:28]
  assign _T_39 = io_Src_A ^ _GEN_0; // @[ALU.scala 60:28]
  assign _GEN_1 = {{63'd0}, io_Src_A}; // @[ALU.scala 61:28]
  assign _T_40 = _GEN_1 << shamt; // @[ALU.scala 61:28]
  assign _T_41 = io_Src_A >> shamt; // @[ALU.scala 62:28]
  assign _T_42 = $signed(io_Src_A); // @[ALU.scala 63:34]
  assign _T_43 = $signed(_T_42) >>> shamt; // @[ALU.scala 63:37]
  assign _T_44 = $unsigned(_T_43); // @[ALU.scala 63:53]
  assign _T_46 = $signed(io_Src_B); // @[ALU.scala 64:54]
  assign _T_47 = $signed(_T_42) < $signed(_T_46); // @[ALU.scala 64:37]
  assign _T_48 = io_Src_A < io_Src_B; // @[ALU.scala 65:28]
  assign _T_49 = 5'h9 == io_ALUOp; // @[Mux.scala 46:19]
  assign _T_50 = _T_49 ? {{31'd0}, _T_48} : io_Src_B; // @[Mux.scala 46:16]
  assign _T_51 = 5'h8 == io_ALUOp; // @[Mux.scala 46:19]
  assign _T_52 = _T_51 ? {{31'd0}, _T_47} : _T_50; // @[Mux.scala 46:16]
  assign _T_53 = 5'h7 == io_ALUOp; // @[Mux.scala 46:19]
  assign _T_54 = _T_53 ? _T_44 : _T_52; // @[Mux.scala 46:16]
  assign _T_55 = 5'h6 == io_ALUOp; // @[Mux.scala 46:19]
  assign _T_56 = _T_55 ? _T_41 : _T_54; // @[Mux.scala 46:16]
  assign _T_57 = 5'h5 == io_ALUOp; // @[Mux.scala 46:19]
  assign _T_58 = _T_57 ? _T_40 : {{63'd0}, _T_56}; // @[Mux.scala 46:16]
  assign _T_59 = 5'h4 == io_ALUOp; // @[Mux.scala 46:19]
  assign _T_60 = _T_59 ? {{63'd0}, _T_39} : _T_58; // @[Mux.scala 46:16]
  assign _T_61 = 5'h3 == io_ALUOp; // @[Mux.scala 46:19]
  assign _T_62 = _T_61 ? {{63'd0}, _T_38} : _T_60; // @[Mux.scala 46:16]
  assign _T_63 = 5'h2 == io_ALUOp; // @[Mux.scala 46:19]
  assign _T_64 = _T_63 ? {{63'd0}, _T_37} : _T_62; // @[Mux.scala 46:16]
  assign _T_65 = 5'h1 == io_ALUOp; // @[Mux.scala 46:19]
  assign _T_66 = _T_65 ? {{63'd0}, _T_36} : _T_64; // @[Mux.scala 46:16]
  assign _T_67 = 5'h0 == io_ALUOp; // @[Mux.scala 46:19]
  assign _T_68 = _T_67 ? {{63'd0}, _T_33} : _T_66; // @[Mux.scala 46:16]
  assign _T_72 = $signed(_T_42) == $signed(_T_46); // @[ALU.scala 69:37]
  assign _T_75 = $signed(_T_42) != $signed(_T_46); // @[ALU.scala 70:37]
  assign _T_81 = $signed(_T_42) >= $signed(_T_46); // @[ALU.scala 72:37]
  assign _T_83 = io_Src_A >= io_Src_B; // @[ALU.scala 74:28]
  assign _T_84 = 5'hf == io_ALUOp; // @[Mux.scala 46:19]
  assign _T_85 = _T_84 ? _T_83 : 1'h0; // @[Mux.scala 46:16]
  assign _T_86 = 5'he == io_ALUOp; // @[Mux.scala 46:19]
  assign _T_87 = _T_86 ? _T_48 : _T_85; // @[Mux.scala 46:16]
  assign _T_88 = 5'hd == io_ALUOp; // @[Mux.scala 46:19]
  assign _T_89 = _T_88 ? _T_81 : _T_87; // @[Mux.scala 46:16]
  assign _T_90 = 5'hc == io_ALUOp; // @[Mux.scala 46:19]
  assign _T_91 = _T_90 ? _T_47 : _T_89; // @[Mux.scala 46:16]
  assign _T_92 = 5'hb == io_ALUOp; // @[Mux.scala 46:19]
  assign _T_93 = _T_92 ? _T_75 : _T_91; // @[Mux.scala 46:16]
  assign _T_94 = 5'ha == io_ALUOp; // @[Mux.scala 46:19]
  assign io_Sum = _T_68[31:0]; // @[ALU.scala 55:10]
  assign io_Conflag = _T_94 ? _T_72 : _T_93; // @[ALU.scala 68:14]
endmodule
