module PC( // @[pc.py:20:Tile.fir@2.2]
  input         clock, // @[rawmodule.py:100:Tile.fir@3.4]
  input         reset, // @[rawmodule.py:101:Tile.fir@4.4]
  input  [31:0] io_next_pc, // @[pc.py:12:Tile.fir@5.4]
  input         io_PC_Write, // @[pc.py:12:Tile.fir@5.4]
  output [31:0] io_pc_out // @[pc.py:12:Tile.fir@5.4]
);
  reg [31:0] pc_reg; // @[pc.py:23:Tile.fir@7.4]
  reg [31:0] _RAND_0;
  assign io_pc_out = pc_reg; // @[pc.py:25:Tile.fir@11.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pc_reg = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      pc_reg <= 32'h0;
    end else begin
      if (io_PC_Write) begin
        pc_reg <= io_next_pc;
      end
    end
  end
endmodule
module InstCache( // @[instcache.py:19:Tile.fir@14.2]
  input         clock, // @[rawmodule.py:100:Tile.fir@15.4]
  input  [31:0] io_addr, // @[instcache.py:12:Tile.fir@17.4]
  output [31:0] io_inst // @[instcache.py:12:Tile.fir@17.4]
);
  reg [7:0] cache [0:1023]; // @[instcache.py:22:Tile.fir@19.4]
  reg [31:0] _RAND_0;
  wire [7:0] cache__T_49_data; // @[instcache.py:22:Tile.fir@19.4]
  wire [9:0] cache__T_49_addr; // @[instcache.py:22:Tile.fir@19.4]
  wire [7:0] cache__T_51_data; // @[instcache.py:22:Tile.fir@19.4]
  wire [9:0] cache__T_51_addr; // @[instcache.py:22:Tile.fir@19.4]
  wire [7:0] cache__T_53_data; // @[instcache.py:22:Tile.fir@19.4]
  wire [9:0] cache__T_53_addr; // @[instcache.py:22:Tile.fir@19.4]
  wire [7:0] cache__T_55_data; // @[instcache.py:22:Tile.fir@19.4]
  wire [9:0] cache__T_55_addr; // @[instcache.py:22:Tile.fir@19.4]
  wire [32:0] _T_50; // @[instcache.py:23:Tile.fir@21.4]
  wire [32:0] _T_52; // @[instcache.py:24:Tile.fir@23.4]
  wire [32:0] _T_54; // @[instcache.py:24:Tile.fir@25.4]
  wire [23:0] _T_57; // @[instcache.py:24:Tile.fir@28.4]
  assign cache__T_49_addr = io_addr[9:0];
  assign cache__T_49_data = cache[cache__T_49_addr]; // @[instcache.py:22:Tile.fir@19.4]
  assign cache__T_51_addr = _T_50[9:0];
  assign cache__T_51_data = cache[cache__T_51_addr]; // @[instcache.py:22:Tile.fir@19.4]
  assign cache__T_53_addr = _T_52[9:0];
  assign cache__T_53_data = cache[cache__T_53_addr]; // @[instcache.py:22:Tile.fir@19.4]
  assign cache__T_55_addr = _T_54[9:0];
  assign cache__T_55_data = cache[cache__T_55_addr]; // @[instcache.py:22:Tile.fir@19.4]
  assign _T_50 = io_addr + 32'h1; // @[instcache.py:23:Tile.fir@21.4]
  assign _T_52 = io_addr + 32'h2; // @[instcache.py:24:Tile.fir@23.4]
  assign _T_54 = io_addr + 32'h3; // @[instcache.py:24:Tile.fir@25.4]
  assign _T_57 = {cache__T_49_data,cache__T_51_data,cache__T_53_data}; // @[instcache.py:24:Tile.fir@28.4]
  assign io_inst = {_T_57,cache__T_55_data}; // @[instcache.py:24:Tile.fir@30.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    cache[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end
endmodule
module Datapath( // @[datapath.py:30:Tile.fir@33.2]
  input  [31:0] io_if_io_pc_out, // @[datapath.py:24:Tile.fir@36.4]
  input  [31:0] io_if_io_pc_recover, // @[datapath.py:24:Tile.fir@36.4]
  input  [31:0] io_if_io_new_addr, // @[datapath.py:24:Tile.fir@36.4]
  output [31:0] io_if_io_next_pc, // @[datapath.py:24:Tile.fir@36.4]
  output [31:0] io_if_io_pc_4, // @[datapath.py:24:Tile.fir@36.4]
  input  [1:0]  io_if_io_PC_Sel // @[datapath.py:24:Tile.fir@36.4]
);
  wire [32:0] _T_71; // @[datapath.py:33:Tile.fir@38.4]
  wire  _T_72; // @[mux.py:72:Tile.fir@40.4]
  wire [31:0] _T_73; // @[datapath.py:38:Tile.fir@41.4]
  wire  _T_74; // @[mux.py:72:Tile.fir@42.4]
  wire [31:0] _T_75; // @[datapath.py:38:Tile.fir@43.4]
  wire  _T_76; // @[mux.py:72:Tile.fir@44.4]
  assign _T_71 = io_if_io_pc_out + 32'h4; // @[datapath.py:33:Tile.fir@38.4]
  assign _T_72 = io_if_io_PC_Sel == 2'h2; // @[mux.py:72:Tile.fir@40.4]
  assign _T_73 = _T_72 ? io_if_io_new_addr : 32'h0; // @[datapath.py:38:Tile.fir@41.4]
  assign _T_74 = io_if_io_PC_Sel == 2'h1; // @[mux.py:72:Tile.fir@42.4]
  assign _T_75 = _T_74 ? io_if_io_pc_recover : _T_73; // @[datapath.py:38:Tile.fir@43.4]
  assign _T_76 = io_if_io_PC_Sel == 2'h0; // @[mux.py:72:Tile.fir@44.4]
  assign io_if_io_next_pc = _T_76 ? io_if_io_pc_4 : _T_75; // @[datapath.py:38:Tile.fir@46.4]
  assign io_if_io_pc_4 = _T_71[31:0]; // @[datapath.py:33:Tile.fir@39.4]
endmodule
module IF_ID_Register( // @[if_id_register.py:28:Tile.fir@49.2]
  input         clock, // @[rawmodule.py:100:Tile.fir@50.4]
  input         reset, // @[rawmodule.py:101:Tile.fir@51.4]
  input  [31:0] io_if_pc, // @[if_id_register.py:11:Tile.fir@52.4]
  input  [31:0] io_if_pc_4, // @[if_id_register.py:11:Tile.fir@52.4]
  input  [31:0] io_if_inst, // @[if_id_register.py:11:Tile.fir@52.4]
  output [31:0] io_id_pc, // @[if_id_register.py:11:Tile.fir@52.4]
  output [31:0] io_id_pc_4, // @[if_id_register.py:11:Tile.fir@52.4]
  output [4:0]  io_id_rs1, // @[if_id_register.py:11:Tile.fir@52.4]
  output [4:0]  io_id_rs2, // @[if_id_register.py:11:Tile.fir@52.4]
  output [31:0] io_id_inst, // @[if_id_register.py:11:Tile.fir@52.4]
  input         io_IF_ID_Write, // @[if_id_register.py:11:Tile.fir@52.4]
  input         io_IF_ID_Flush // @[if_id_register.py:11:Tile.fir@52.4]
);
  reg [31:0] pc; // @[if_id_register.py:31:Tile.fir@54.4]
  reg [31:0] _RAND_0;
  reg [31:0] pc_4; // @[if_id_register.py:32:Tile.fir@55.4]
  reg [31:0] _RAND_1;
  reg [31:0] inst; // @[if_id_register.py:33:Tile.fir@56.4]
  reg [31:0] _RAND_2;
  assign io_id_pc = pc; // @[if_id_register.py:42:Tile.fir@72.4]
  assign io_id_pc_4 = pc_4; // @[if_id_register.py:43:Tile.fir@73.4]
  assign io_id_rs1 = inst[19:15]; // @[if_id_register.py:45:Tile.fir@76.4]
  assign io_id_rs2 = inst[24:20]; // @[if_id_register.py:46:Tile.fir@78.4]
  assign io_id_inst = inst; // @[if_id_register.py:44:Tile.fir@74.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pc = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  pc_4 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  inst = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      pc <= 32'h0;
    end else begin
      if (io_IF_ID_Flush) begin
        pc <= 32'h0;
      end else begin
        if (io_IF_ID_Write) begin
          pc <= io_if_pc;
        end
      end
    end
    if (reset) begin
      pc_4 <= 32'h0;
    end else begin
      if (io_IF_ID_Flush) begin
        pc_4 <= 32'h0;
      end else begin
        if (io_IF_ID_Write) begin
          pc_4 <= io_if_pc_4;
        end
      end
    end
    if (reset) begin
      inst <= 32'h0;
    end else begin
      if (io_IF_ID_Flush) begin
        inst <= 32'h0;
      end else begin
        if (io_IF_ID_Write) begin
          inst <= io_if_inst;
        end
      end
    end
  end
endmodule
module RegFile( // @[regfile.py:24:Tile.fir@81.2]
  input         clock, // @[rawmodule.py:100:Tile.fir@82.4]
  input  [4:0]  io_rs1, // @[regfile.py:11:Tile.fir@84.4]
  input  [4:0]  io_rs2, // @[regfile.py:11:Tile.fir@84.4]
  input  [4:0]  io_rd, // @[regfile.py:11:Tile.fir@84.4]
  input  [31:0] io_wdata, // @[regfile.py:11:Tile.fir@84.4]
  output [31:0] io_rs1_out, // @[regfile.py:11:Tile.fir@84.4]
  output [31:0] io_rs2_out, // @[regfile.py:11:Tile.fir@84.4]
  input         io_Reg_Write // @[regfile.py:11:Tile.fir@84.4]
);
  reg [31:0] regfile [0:31]; // @[regfile.py:27:Tile.fir@86.4]
  reg [31:0] _RAND_0;
  wire [31:0] regfile__T_127_data; // @[regfile.py:27:Tile.fir@86.4]
  wire [4:0] regfile__T_127_addr; // @[regfile.py:27:Tile.fir@86.4]
  wire [31:0] regfile__T_129_data; // @[regfile.py:27:Tile.fir@86.4]
  wire [4:0] regfile__T_129_addr; // @[regfile.py:27:Tile.fir@86.4]
  wire [31:0] regfile__T_134_data; // @[regfile.py:27:Tile.fir@86.4]
  wire [4:0] regfile__T_134_addr; // @[regfile.py:27:Tile.fir@86.4]
  wire [31:0] regfile__T_136_data; // @[regfile.py:27:Tile.fir@86.4]
  wire [4:0] regfile__T_136_addr; // @[regfile.py:27:Tile.fir@86.4]
  wire  regfile__T_136_mask; // @[regfile.py:27:Tile.fir@86.4]
  wire  regfile__T_136_en; // @[regfile.py:27:Tile.fir@86.4]
  wire  _T_122; // @[regfile.py:30:Tile.fir@88.4]
  wire  _T_123; // @[regfile.py:30:Tile.fir@89.4]
  wire  _T_125; // @[regfile.py:31:Tile.fir@91.4]
  wire  _T_126; // @[regfile.py:31:Tile.fir@92.4]
  wire  _T_132; // @[regfile.py:36:Tile.fir@100.4]
  wire [31:0] _T_133; // @[regfile.py:36:Tile.fir@101.4]
  assign regfile__T_127_addr = io_rs1;
  assign regfile__T_127_data = regfile[regfile__T_127_addr]; // @[regfile.py:27:Tile.fir@86.4]
  assign regfile__T_129_addr = io_rs2;
  assign regfile__T_129_data = regfile[regfile__T_129_addr]; // @[regfile.py:27:Tile.fir@86.4]
  assign regfile__T_134_addr = io_rd;
  assign regfile__T_134_data = regfile[regfile__T_134_addr]; // @[regfile.py:27:Tile.fir@86.4]
  assign regfile__T_136_data = io_Reg_Write ? _T_133 : regfile__T_134_data;
  assign regfile__T_136_addr = io_rd;
  assign regfile__T_136_mask = 1'h1;
  assign regfile__T_136_en = 1'h1;
  assign _T_122 = io_rs1 == io_rd; // @[regfile.py:30:Tile.fir@88.4]
  assign _T_123 = io_Reg_Write & _T_122; // @[regfile.py:30:Tile.fir@89.4]
  assign _T_125 = io_rs2 == io_rd; // @[regfile.py:31:Tile.fir@91.4]
  assign _T_126 = io_Reg_Write & _T_125; // @[regfile.py:31:Tile.fir@92.4]
  assign _T_132 = io_rd == 5'h0; // @[regfile.py:36:Tile.fir@100.4]
  assign _T_133 = _T_132 ? 32'h0 : io_wdata; // @[regfile.py:36:Tile.fir@101.4]
  assign io_rs1_out = _T_123 ? io_wdata : regfile__T_127_data; // @[regfile.py:33:Tile.fir@95.4]
  assign io_rs2_out = _T_126 ? io_wdata : regfile__T_129_data; // @[regfile.py:34:Tile.fir@98.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    regfile[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if(regfile__T_136_en & regfile__T_136_mask) begin
      regfile[regfile__T_136_addr] <= regfile__T_136_data; // @[regfile.py:27:Tile.fir@86.4]
    end
  end
endmodule
module ImmGen( // @[immgen.py:20:Tile.fir@108.2]
  input  [31:0] io_inst, // @[immgen.py:11:Tile.fir@111.4]
  output [31:0] io_imm, // @[immgen.py:11:Tile.fir@111.4]
  input  [2:0]  io_Imm_Sel // @[immgen.py:11:Tile.fir@111.4]
);
  wire [11:0] _T_145; // @[immgen.py:24:Tile.fir@114.4]
  wire [11:0] _T_146; // @[immgen.py:24:Tile.fir@115.4]
  wire [6:0] _T_147; // @[immgen.py:25:Tile.fir@116.4]
  wire [4:0] _T_148; // @[immgen.py:25:Tile.fir@117.4]
  wire [11:0] _T_149; // @[immgen.py:25:Tile.fir@118.4]
  wire [11:0] _T_150; // @[immgen.py:25:Tile.fir@119.4]
  wire  _T_151; // @[immgen.py:26:Tile.fir@120.4]
  wire  _T_152; // @[immgen.py:26:Tile.fir@121.4]
  wire [5:0] _T_153; // @[immgen.py:26:Tile.fir@123.4]
  wire [3:0] _T_154; // @[immgen.py:26:Tile.fir@125.4]
  wire [12:0] _T_158; // @[immgen.py:26:Tile.fir@127.4]
  wire [12:0] _T_159; // @[immgen.py:26:Tile.fir@128.4]
  wire [19:0] _T_160; // @[immgen.py:27:Tile.fir@129.4]
  wire [31:0] _T_161; // @[immgen.py:27:Tile.fir@130.4]
  wire [31:0] _T_162; // @[immgen.py:27:Tile.fir@131.4]
  wire [7:0] _T_164; // @[immgen.py:28:Tile.fir@133.4]
  wire  _T_165; // @[immgen.py:28:Tile.fir@135.4]
  wire [9:0] _T_166; // @[immgen.py:28:Tile.fir@137.4]
  wire [20:0] _T_170; // @[immgen.py:28:Tile.fir@139.4]
  wire [20:0] _T_171; // @[immgen.py:28:Tile.fir@140.4]
  wire  _T_172; // @[mux.py:72:Tile.fir@141.4]
  wire [31:0] _T_173; // @[immgen.py:36:Tile.fir@142.4]
  wire  _T_174; // @[mux.py:72:Tile.fir@143.4]
  wire [31:0] _T_175; // @[immgen.py:36:Tile.fir@144.4]
  wire  _T_176; // @[mux.py:72:Tile.fir@145.4]
  wire [31:0] _T_177; // @[immgen.py:36:Tile.fir@146.4]
  wire  _T_178; // @[mux.py:72:Tile.fir@147.4]
  wire [31:0] _T_179; // @[immgen.py:36:Tile.fir@148.4]
  wire  _T_180; // @[mux.py:72:Tile.fir@149.4]
  wire [31:0] _T_181; // @[immgen.py:36:Tile.fir@150.4]
  wire  _T_182; // @[mux.py:72:Tile.fir@151.4]
  wire [31:0] _T_183; // @[immgen.py:36:Tile.fir@152.4]
  assign _T_145 = io_inst[31:20]; // @[immgen.py:24:Tile.fir@114.4]
  assign _T_146 = $signed(_T_145); // @[immgen.py:24:Tile.fir@115.4]
  assign _T_147 = io_inst[31:25]; // @[immgen.py:25:Tile.fir@116.4]
  assign _T_148 = io_inst[11:7]; // @[immgen.py:25:Tile.fir@117.4]
  assign _T_149 = {_T_147,_T_148}; // @[immgen.py:25:Tile.fir@118.4]
  assign _T_150 = $signed(_T_149); // @[immgen.py:25:Tile.fir@119.4]
  assign _T_151 = io_inst[31]; // @[immgen.py:26:Tile.fir@120.4]
  assign _T_152 = io_inst[7]; // @[immgen.py:26:Tile.fir@121.4]
  assign _T_153 = io_inst[30:25]; // @[immgen.py:26:Tile.fir@123.4]
  assign _T_154 = io_inst[11:8]; // @[immgen.py:26:Tile.fir@125.4]
  assign _T_158 = {_T_151,_T_152,_T_153,_T_154,1'h0}; // @[immgen.py:26:Tile.fir@127.4]
  assign _T_159 = $signed(_T_158); // @[immgen.py:26:Tile.fir@128.4]
  assign _T_160 = io_inst[31:12]; // @[immgen.py:27:Tile.fir@129.4]
  assign _T_161 = {_T_160,12'h0}; // @[immgen.py:27:Tile.fir@130.4]
  assign _T_162 = $signed(_T_161); // @[immgen.py:27:Tile.fir@131.4]
  assign _T_164 = io_inst[19:12]; // @[immgen.py:28:Tile.fir@133.4]
  assign _T_165 = io_inst[20]; // @[immgen.py:28:Tile.fir@135.4]
  assign _T_166 = io_inst[30:21]; // @[immgen.py:28:Tile.fir@137.4]
  assign _T_170 = {_T_151,_T_164,_T_165,_T_166,1'h0}; // @[immgen.py:28:Tile.fir@139.4]
  assign _T_171 = $signed(_T_170); // @[immgen.py:28:Tile.fir@140.4]
  assign _T_172 = io_Imm_Sel == 3'h6; // @[mux.py:72:Tile.fir@141.4]
  assign _T_173 = _T_172 ? $signed({{11{_T_171[20]}},_T_171}) : $signed(32'sh0); // @[immgen.py:36:Tile.fir@142.4]
  assign _T_174 = io_Imm_Sel == 3'h5; // @[mux.py:72:Tile.fir@143.4]
  assign _T_175 = _T_174 ? $signed(_T_162) : $signed(_T_173); // @[immgen.py:36:Tile.fir@144.4]
  assign _T_176 = io_Imm_Sel == 3'h4; // @[mux.py:72:Tile.fir@145.4]
  assign _T_177 = _T_176 ? $signed({{19{_T_159[12]}},_T_159}) : $signed(_T_175); // @[immgen.py:36:Tile.fir@146.4]
  assign _T_178 = io_Imm_Sel == 3'h3; // @[mux.py:72:Tile.fir@147.4]
  assign _T_179 = _T_178 ? $signed({{20{_T_150[11]}},_T_150}) : $signed(_T_177); // @[immgen.py:36:Tile.fir@148.4]
  assign _T_180 = io_Imm_Sel == 3'h2; // @[mux.py:72:Tile.fir@149.4]
  assign _T_181 = _T_180 ? $signed({{20{_T_146[11]}},_T_146}) : $signed(_T_179); // @[immgen.py:36:Tile.fir@150.4]
  assign _T_182 = io_Imm_Sel == 3'h1; // @[mux.py:72:Tile.fir@151.4]
  assign _T_183 = _T_182 ? $signed(32'sh0) : $signed(_T_181); // @[immgen.py:36:Tile.fir@152.4]
  assign io_imm = $unsigned(_T_183); // @[immgen.py:36:Tile.fir@154.4]
endmodule
module Control( // @[control.py:86:Tile.fir@157.2]
  input  [31:0] io_inst, // @[control.py:68:Tile.fir@160.4]
  output        io_Reg_Write, // @[control.py:68:Tile.fir@160.4]
  output [2:0]  io_Imm_Sel, // @[control.py:68:Tile.fir@160.4]
  output        io_ALU_Src, // @[control.py:68:Tile.fir@160.4]
  output [4:0]  io_ALUOp, // @[control.py:68:Tile.fir@160.4]
  output        io_Branch, // @[control.py:68:Tile.fir@160.4]
  output        io_Branch_Src, // @[control.py:68:Tile.fir@160.4]
  output        io_Mem_Read, // @[control.py:68:Tile.fir@160.4]
  output        io_Mem_Write, // @[control.py:68:Tile.fir@160.4]
  output [1:0]  io_Data_Size, // @[control.py:68:Tile.fir@160.4]
  output        io_Load_Type, // @[control.py:68:Tile.fir@160.4]
  output [2:0]  io_Mem_to_Reg, // @[control.py:68:Tile.fir@160.4]
  output        io_Jump_Type // @[control.py:68:Tile.fir@160.4]
);
  wire [31:0] _T_202; // @[listlookup.py:52:Tile.fir@162.4]
  wire  _T_203; // @[listlookup.py:52:Tile.fir@163.4]
  wire  _T_205; // @[listlookup.py:52:Tile.fir@165.4]
  wire  _T_207; // @[listlookup.py:52:Tile.fir@167.4]
  wire  _T_209; // @[listlookup.py:52:Tile.fir@169.4]
  wire  _T_211; // @[listlookup.py:52:Tile.fir@171.4]
  wire [31:0] _T_212; // @[listlookup.py:52:Tile.fir@172.4]
  wire  _T_213; // @[listlookup.py:52:Tile.fir@173.4]
  wire  _T_215; // @[listlookup.py:52:Tile.fir@175.4]
  wire  _T_217; // @[listlookup.py:52:Tile.fir@177.4]
  wire  _T_219; // @[listlookup.py:52:Tile.fir@179.4]
  wire  _T_221; // @[listlookup.py:52:Tile.fir@181.4]
  wire  _T_223; // @[listlookup.py:52:Tile.fir@183.4]
  wire  _T_225; // @[listlookup.py:52:Tile.fir@185.4]
  wire  _T_227; // @[listlookup.py:52:Tile.fir@187.4]
  wire  _T_229; // @[listlookup.py:52:Tile.fir@189.4]
  wire  _T_231; // @[listlookup.py:52:Tile.fir@191.4]
  wire  _T_233; // @[listlookup.py:52:Tile.fir@193.4]
  wire  _T_235; // @[listlookup.py:52:Tile.fir@195.4]
  wire  _T_237; // @[listlookup.py:52:Tile.fir@197.4]
  wire  _T_239; // @[listlookup.py:52:Tile.fir@199.4]
  wire  _T_241; // @[listlookup.py:52:Tile.fir@201.4]
  wire  _T_243; // @[listlookup.py:52:Tile.fir@203.4]
  wire  _T_245; // @[listlookup.py:52:Tile.fir@205.4]
  wire  _T_247; // @[listlookup.py:52:Tile.fir@207.4]
  wire  _T_249; // @[listlookup.py:52:Tile.fir@209.4]
  wire  _T_251; // @[listlookup.py:52:Tile.fir@211.4]
  wire  _T_253; // @[listlookup.py:52:Tile.fir@213.4]
  wire  _T_255; // @[listlookup.py:52:Tile.fir@215.4]
  wire  _T_257; // @[listlookup.py:52:Tile.fir@217.4]
  wire  _T_259; // @[listlookup.py:52:Tile.fir@219.4]
  wire  _T_261; // @[listlookup.py:52:Tile.fir@221.4]
  wire  _T_263; // @[listlookup.py:52:Tile.fir@223.4]
  wire  _T_265; // @[listlookup.py:52:Tile.fir@225.4]
  wire  _T_267; // @[listlookup.py:52:Tile.fir@227.4]
  wire [31:0] _T_268; // @[listlookup.py:52:Tile.fir@228.4]
  wire  _T_269; // @[listlookup.py:52:Tile.fir@229.4]
  wire  _T_271; // @[listlookup.py:52:Tile.fir@231.4]
  wire  _T_273; // @[listlookup.py:52:Tile.fir@233.4]
  wire  _T_275; // @[listlookup.py:52:Tile.fir@235.4]
  wire  _T_280; // @[control.py:89:Tile.fir@240.4]
  wire  _T_281; // @[control.py:89:Tile.fir@241.4]
  wire  _T_282; // @[control.py:89:Tile.fir@242.4]
  wire  _T_283; // @[control.py:89:Tile.fir@243.4]
  wire  _T_284; // @[control.py:89:Tile.fir@244.4]
  wire  _T_285; // @[control.py:89:Tile.fir@245.4]
  wire  _T_286; // @[control.py:89:Tile.fir@246.4]
  wire  _T_287; // @[control.py:89:Tile.fir@247.4]
  wire  _T_288; // @[control.py:89:Tile.fir@248.4]
  wire  _T_289; // @[control.py:89:Tile.fir@249.4]
  wire  _T_290; // @[control.py:89:Tile.fir@250.4]
  wire  _T_291; // @[control.py:89:Tile.fir@251.4]
  wire  _T_292; // @[control.py:89:Tile.fir@252.4]
  wire  _T_293; // @[control.py:89:Tile.fir@253.4]
  wire  _T_294; // @[control.py:89:Tile.fir@254.4]
  wire  _T_295; // @[control.py:89:Tile.fir@255.4]
  wire  _T_296; // @[control.py:89:Tile.fir@256.4]
  wire  _T_297; // @[control.py:89:Tile.fir@257.4]
  wire  _T_298; // @[control.py:89:Tile.fir@258.4]
  wire  _T_299; // @[control.py:89:Tile.fir@259.4]
  wire  _T_300; // @[control.py:89:Tile.fir@260.4]
  wire  _T_301; // @[control.py:89:Tile.fir@261.4]
  wire  _T_302; // @[control.py:89:Tile.fir@262.4]
  wire  _T_303; // @[control.py:89:Tile.fir@263.4]
  wire  _T_304; // @[control.py:89:Tile.fir@264.4]
  wire  _T_305; // @[control.py:89:Tile.fir@265.4]
  wire  _T_306; // @[control.py:89:Tile.fir@266.4]
  wire  _T_307; // @[control.py:89:Tile.fir@267.4]
  wire  _T_308; // @[control.py:89:Tile.fir@268.4]
  wire  _T_309; // @[control.py:89:Tile.fir@269.4]
  wire  _T_310; // @[control.py:89:Tile.fir@270.4]
  wire  _T_311; // @[control.py:89:Tile.fir@271.4]
  wire  _T_312; // @[control.py:89:Tile.fir@272.4]
  wire  _T_313; // @[control.py:89:Tile.fir@273.4]
  wire  _T_314; // @[control.py:89:Tile.fir@274.4]
  wire [2:0] _T_317; // @[control.py:89:Tile.fir@277.4]
  wire [2:0] _T_318; // @[control.py:89:Tile.fir@278.4]
  wire [2:0] _T_319; // @[control.py:89:Tile.fir@279.4]
  wire [2:0] _T_320; // @[control.py:89:Tile.fir@280.4]
  wire [2:0] _T_321; // @[control.py:89:Tile.fir@281.4]
  wire [2:0] _T_322; // @[control.py:89:Tile.fir@282.4]
  wire [2:0] _T_323; // @[control.py:89:Tile.fir@283.4]
  wire [2:0] _T_324; // @[control.py:89:Tile.fir@284.4]
  wire [2:0] _T_325; // @[control.py:89:Tile.fir@285.4]
  wire [2:0] _T_326; // @[control.py:89:Tile.fir@286.4]
  wire [2:0] _T_327; // @[control.py:89:Tile.fir@287.4]
  wire [2:0] _T_328; // @[control.py:89:Tile.fir@288.4]
  wire [2:0] _T_329; // @[control.py:89:Tile.fir@289.4]
  wire [2:0] _T_330; // @[control.py:89:Tile.fir@290.4]
  wire [2:0] _T_331; // @[control.py:89:Tile.fir@291.4]
  wire [2:0] _T_332; // @[control.py:89:Tile.fir@292.4]
  wire [2:0] _T_333; // @[control.py:89:Tile.fir@293.4]
  wire [2:0] _T_334; // @[control.py:89:Tile.fir@294.4]
  wire [2:0] _T_335; // @[control.py:89:Tile.fir@295.4]
  wire [2:0] _T_336; // @[control.py:89:Tile.fir@296.4]
  wire [2:0] _T_337; // @[control.py:89:Tile.fir@297.4]
  wire [2:0] _T_338; // @[control.py:89:Tile.fir@298.4]
  wire [2:0] _T_339; // @[control.py:89:Tile.fir@299.4]
  wire [2:0] _T_340; // @[control.py:89:Tile.fir@300.4]
  wire [2:0] _T_341; // @[control.py:89:Tile.fir@301.4]
  wire [2:0] _T_342; // @[control.py:89:Tile.fir@302.4]
  wire [2:0] _T_343; // @[control.py:89:Tile.fir@303.4]
  wire [2:0] _T_344; // @[control.py:89:Tile.fir@304.4]
  wire [2:0] _T_345; // @[control.py:89:Tile.fir@305.4]
  wire [2:0] _T_346; // @[control.py:89:Tile.fir@306.4]
  wire [2:0] _T_347; // @[control.py:89:Tile.fir@307.4]
  wire [2:0] _T_348; // @[control.py:89:Tile.fir@308.4]
  wire [2:0] _T_349; // @[control.py:89:Tile.fir@309.4]
  wire [2:0] _T_350; // @[control.py:89:Tile.fir@310.4]
  wire [2:0] _T_351; // @[control.py:89:Tile.fir@311.4]
  wire [2:0] _T_352; // @[control.py:89:Tile.fir@312.4]
  wire  _T_366; // @[control.py:89:Tile.fir@326.4]
  wire  _T_367; // @[control.py:89:Tile.fir@327.4]
  wire  _T_368; // @[control.py:89:Tile.fir@328.4]
  wire  _T_369; // @[control.py:89:Tile.fir@329.4]
  wire  _T_370; // @[control.py:89:Tile.fir@330.4]
  wire  _T_371; // @[control.py:89:Tile.fir@331.4]
  wire  _T_372; // @[control.py:89:Tile.fir@332.4]
  wire  _T_373; // @[control.py:89:Tile.fir@333.4]
  wire  _T_374; // @[control.py:89:Tile.fir@334.4]
  wire  _T_375; // @[control.py:89:Tile.fir@335.4]
  wire  _T_376; // @[control.py:89:Tile.fir@336.4]
  wire  _T_377; // @[control.py:89:Tile.fir@337.4]
  wire  _T_378; // @[control.py:89:Tile.fir@338.4]
  wire  _T_379; // @[control.py:89:Tile.fir@339.4]
  wire  _T_380; // @[control.py:89:Tile.fir@340.4]
  wire  _T_381; // @[control.py:89:Tile.fir@341.4]
  wire  _T_382; // @[control.py:89:Tile.fir@342.4]
  wire  _T_383; // @[control.py:89:Tile.fir@343.4]
  wire  _T_384; // @[control.py:89:Tile.fir@344.4]
  wire  _T_385; // @[control.py:89:Tile.fir@345.4]
  wire  _T_386; // @[control.py:89:Tile.fir@346.4]
  wire  _T_387; // @[control.py:89:Tile.fir@347.4]
  wire  _T_388; // @[control.py:89:Tile.fir@348.4]
  wire  _T_389; // @[control.py:89:Tile.fir@349.4]
  wire  _T_390; // @[control.py:89:Tile.fir@350.4]
  wire [4:0] _T_393; // @[control.py:89:Tile.fir@353.4]
  wire [4:0] _T_394; // @[control.py:89:Tile.fir@354.4]
  wire [4:0] _T_395; // @[control.py:89:Tile.fir@355.4]
  wire [4:0] _T_396; // @[control.py:89:Tile.fir@356.4]
  wire [4:0] _T_397; // @[control.py:89:Tile.fir@357.4]
  wire [4:0] _T_398; // @[control.py:89:Tile.fir@358.4]
  wire [4:0] _T_399; // @[control.py:89:Tile.fir@359.4]
  wire [4:0] _T_400; // @[control.py:89:Tile.fir@360.4]
  wire [4:0] _T_401; // @[control.py:89:Tile.fir@361.4]
  wire [4:0] _T_402; // @[control.py:89:Tile.fir@362.4]
  wire [4:0] _T_403; // @[control.py:89:Tile.fir@363.4]
  wire [4:0] _T_404; // @[control.py:89:Tile.fir@364.4]
  wire [4:0] _T_405; // @[control.py:89:Tile.fir@365.4]
  wire [4:0] _T_406; // @[control.py:89:Tile.fir@366.4]
  wire [4:0] _T_407; // @[control.py:89:Tile.fir@367.4]
  wire [4:0] _T_408; // @[control.py:89:Tile.fir@368.4]
  wire [4:0] _T_409; // @[control.py:89:Tile.fir@369.4]
  wire [4:0] _T_410; // @[control.py:89:Tile.fir@370.4]
  wire [4:0] _T_411; // @[control.py:89:Tile.fir@371.4]
  wire [4:0] _T_412; // @[control.py:89:Tile.fir@372.4]
  wire [4:0] _T_413; // @[control.py:89:Tile.fir@373.4]
  wire [4:0] _T_414; // @[control.py:89:Tile.fir@374.4]
  wire [4:0] _T_415; // @[control.py:89:Tile.fir@375.4]
  wire [4:0] _T_416; // @[control.py:89:Tile.fir@376.4]
  wire [4:0] _T_417; // @[control.py:89:Tile.fir@377.4]
  wire [4:0] _T_418; // @[control.py:89:Tile.fir@378.4]
  wire [4:0] _T_419; // @[control.py:89:Tile.fir@379.4]
  wire [4:0] _T_420; // @[control.py:89:Tile.fir@380.4]
  wire [4:0] _T_421; // @[control.py:89:Tile.fir@381.4]
  wire [4:0] _T_422; // @[control.py:89:Tile.fir@382.4]
  wire [4:0] _T_423; // @[control.py:89:Tile.fir@383.4]
  wire [4:0] _T_424; // @[control.py:89:Tile.fir@384.4]
  wire [4:0] _T_425; // @[control.py:89:Tile.fir@385.4]
  wire [4:0] _T_426; // @[control.py:89:Tile.fir@386.4]
  wire [4:0] _T_427; // @[control.py:89:Tile.fir@387.4]
  wire [4:0] _T_428; // @[control.py:89:Tile.fir@388.4]
  wire  _T_434; // @[control.py:89:Tile.fir@394.4]
  wire  _T_435; // @[control.py:89:Tile.fir@395.4]
  wire  _T_436; // @[control.py:89:Tile.fir@396.4]
  wire  _T_437; // @[control.py:89:Tile.fir@397.4]
  wire  _T_438; // @[control.py:89:Tile.fir@398.4]
  wire  _T_439; // @[control.py:89:Tile.fir@399.4]
  wire  _T_440; // @[control.py:89:Tile.fir@400.4]
  wire  _T_441; // @[control.py:89:Tile.fir@401.4]
  wire  _T_442; // @[control.py:89:Tile.fir@402.4]
  wire  _T_443; // @[control.py:89:Tile.fir@403.4]
  wire  _T_444; // @[control.py:89:Tile.fir@404.4]
  wire  _T_445; // @[control.py:89:Tile.fir@405.4]
  wire  _T_446; // @[control.py:89:Tile.fir@406.4]
  wire  _T_447; // @[control.py:89:Tile.fir@407.4]
  wire  _T_448; // @[control.py:89:Tile.fir@408.4]
  wire  _T_449; // @[control.py:89:Tile.fir@409.4]
  wire  _T_450; // @[control.py:89:Tile.fir@410.4]
  wire  _T_451; // @[control.py:89:Tile.fir@411.4]
  wire  _T_452; // @[control.py:89:Tile.fir@412.4]
  wire  _T_453; // @[control.py:89:Tile.fir@413.4]
  wire  _T_454; // @[control.py:89:Tile.fir@414.4]
  wire  _T_455; // @[control.py:89:Tile.fir@415.4]
  wire  _T_456; // @[control.py:89:Tile.fir@416.4]
  wire  _T_457; // @[control.py:89:Tile.fir@417.4]
  wire  _T_458; // @[control.py:89:Tile.fir@418.4]
  wire  _T_459; // @[control.py:89:Tile.fir@419.4]
  wire  _T_460; // @[control.py:89:Tile.fir@420.4]
  wire  _T_461; // @[control.py:89:Tile.fir@421.4]
  wire  _T_462; // @[control.py:89:Tile.fir@422.4]
  wire  _T_463; // @[control.py:89:Tile.fir@423.4]
  wire  _T_464; // @[control.py:89:Tile.fir@424.4]
  wire  _T_465; // @[control.py:89:Tile.fir@425.4]
  wire  _T_466; // @[control.py:89:Tile.fir@426.4]
  wire  _T_472; // @[control.py:89:Tile.fir@432.4]
  wire  _T_473; // @[control.py:89:Tile.fir@433.4]
  wire  _T_474; // @[control.py:89:Tile.fir@434.4]
  wire  _T_475; // @[control.py:89:Tile.fir@435.4]
  wire  _T_476; // @[control.py:89:Tile.fir@436.4]
  wire  _T_477; // @[control.py:89:Tile.fir@437.4]
  wire  _T_478; // @[control.py:89:Tile.fir@438.4]
  wire  _T_479; // @[control.py:89:Tile.fir@439.4]
  wire  _T_480; // @[control.py:89:Tile.fir@440.4]
  wire  _T_481; // @[control.py:89:Tile.fir@441.4]
  wire  _T_482; // @[control.py:89:Tile.fir@442.4]
  wire  _T_483; // @[control.py:89:Tile.fir@443.4]
  wire  _T_484; // @[control.py:89:Tile.fir@444.4]
  wire  _T_485; // @[control.py:89:Tile.fir@445.4]
  wire  _T_486; // @[control.py:89:Tile.fir@446.4]
  wire  _T_487; // @[control.py:89:Tile.fir@447.4]
  wire  _T_488; // @[control.py:89:Tile.fir@448.4]
  wire  _T_489; // @[control.py:89:Tile.fir@449.4]
  wire  _T_490; // @[control.py:89:Tile.fir@450.4]
  wire  _T_491; // @[control.py:89:Tile.fir@451.4]
  wire  _T_492; // @[control.py:89:Tile.fir@452.4]
  wire  _T_493; // @[control.py:89:Tile.fir@453.4]
  wire  _T_494; // @[control.py:89:Tile.fir@454.4]
  wire  _T_495; // @[control.py:89:Tile.fir@455.4]
  wire  _T_496; // @[control.py:89:Tile.fir@456.4]
  wire  _T_497; // @[control.py:89:Tile.fir@457.4]
  wire  _T_498; // @[control.py:89:Tile.fir@458.4]
  wire  _T_499; // @[control.py:89:Tile.fir@459.4]
  wire  _T_500; // @[control.py:89:Tile.fir@460.4]
  wire  _T_501; // @[control.py:89:Tile.fir@461.4]
  wire  _T_502; // @[control.py:89:Tile.fir@462.4]
  wire  _T_503; // @[control.py:89:Tile.fir@463.4]
  wire  _T_504; // @[control.py:89:Tile.fir@464.4]
  wire  _T_521; // @[control.py:89:Tile.fir@481.4]
  wire  _T_522; // @[control.py:89:Tile.fir@482.4]
  wire  _T_523; // @[control.py:89:Tile.fir@483.4]
  wire  _T_524; // @[control.py:89:Tile.fir@484.4]
  wire  _T_525; // @[control.py:89:Tile.fir@485.4]
  wire  _T_526; // @[control.py:89:Tile.fir@486.4]
  wire  _T_527; // @[control.py:89:Tile.fir@487.4]
  wire  _T_528; // @[control.py:89:Tile.fir@488.4]
  wire  _T_529; // @[control.py:89:Tile.fir@489.4]
  wire  _T_530; // @[control.py:89:Tile.fir@490.4]
  wire  _T_531; // @[control.py:89:Tile.fir@491.4]
  wire  _T_532; // @[control.py:89:Tile.fir@492.4]
  wire  _T_533; // @[control.py:89:Tile.fir@493.4]
  wire  _T_534; // @[control.py:89:Tile.fir@494.4]
  wire  _T_535; // @[control.py:89:Tile.fir@495.4]
  wire  _T_536; // @[control.py:89:Tile.fir@496.4]
  wire  _T_537; // @[control.py:89:Tile.fir@497.4]
  wire  _T_538; // @[control.py:89:Tile.fir@498.4]
  wire  _T_539; // @[control.py:89:Tile.fir@499.4]
  wire  _T_540; // @[control.py:89:Tile.fir@500.4]
  wire  _T_541; // @[control.py:89:Tile.fir@501.4]
  wire  _T_542; // @[control.py:89:Tile.fir@502.4]
  wire  _T_558; // @[control.py:89:Tile.fir@518.4]
  wire  _T_559; // @[control.py:89:Tile.fir@519.4]
  wire  _T_560; // @[control.py:89:Tile.fir@520.4]
  wire  _T_561; // @[control.py:89:Tile.fir@521.4]
  wire  _T_562; // @[control.py:89:Tile.fir@522.4]
  wire  _T_563; // @[control.py:89:Tile.fir@523.4]
  wire  _T_564; // @[control.py:89:Tile.fir@524.4]
  wire  _T_565; // @[control.py:89:Tile.fir@525.4]
  wire  _T_566; // @[control.py:89:Tile.fir@526.4]
  wire  _T_567; // @[control.py:89:Tile.fir@527.4]
  wire  _T_568; // @[control.py:89:Tile.fir@528.4]
  wire  _T_569; // @[control.py:89:Tile.fir@529.4]
  wire  _T_570; // @[control.py:89:Tile.fir@530.4]
  wire  _T_571; // @[control.py:89:Tile.fir@531.4]
  wire  _T_572; // @[control.py:89:Tile.fir@532.4]
  wire  _T_573; // @[control.py:89:Tile.fir@533.4]
  wire  _T_574; // @[control.py:89:Tile.fir@534.4]
  wire  _T_575; // @[control.py:89:Tile.fir@535.4]
  wire  _T_576; // @[control.py:89:Tile.fir@536.4]
  wire  _T_577; // @[control.py:89:Tile.fir@537.4]
  wire  _T_578; // @[control.py:89:Tile.fir@538.4]
  wire  _T_579; // @[control.py:89:Tile.fir@539.4]
  wire  _T_580; // @[control.py:89:Tile.fir@540.4]
  wire [1:0] _T_593; // @[control.py:89:Tile.fir@553.4]
  wire [1:0] _T_594; // @[control.py:89:Tile.fir@554.4]
  wire [1:0] _T_595; // @[control.py:89:Tile.fir@555.4]
  wire [1:0] _T_596; // @[control.py:89:Tile.fir@556.4]
  wire [1:0] _T_597; // @[control.py:89:Tile.fir@557.4]
  wire [1:0] _T_598; // @[control.py:89:Tile.fir@558.4]
  wire [1:0] _T_599; // @[control.py:89:Tile.fir@559.4]
  wire [1:0] _T_600; // @[control.py:89:Tile.fir@560.4]
  wire [1:0] _T_601; // @[control.py:89:Tile.fir@561.4]
  wire [1:0] _T_602; // @[control.py:89:Tile.fir@562.4]
  wire [1:0] _T_603; // @[control.py:89:Tile.fir@563.4]
  wire [1:0] _T_604; // @[control.py:89:Tile.fir@564.4]
  wire [1:0] _T_605; // @[control.py:89:Tile.fir@565.4]
  wire [1:0] _T_606; // @[control.py:89:Tile.fir@566.4]
  wire [1:0] _T_607; // @[control.py:89:Tile.fir@567.4]
  wire [1:0] _T_608; // @[control.py:89:Tile.fir@568.4]
  wire [1:0] _T_609; // @[control.py:89:Tile.fir@569.4]
  wire [1:0] _T_610; // @[control.py:89:Tile.fir@570.4]
  wire [1:0] _T_611; // @[control.py:89:Tile.fir@571.4]
  wire [1:0] _T_612; // @[control.py:89:Tile.fir@572.4]
  wire [1:0] _T_613; // @[control.py:89:Tile.fir@573.4]
  wire [1:0] _T_614; // @[control.py:89:Tile.fir@574.4]
  wire [1:0] _T_615; // @[control.py:89:Tile.fir@575.4]
  wire [1:0] _T_616; // @[control.py:89:Tile.fir@576.4]
  wire [1:0] _T_617; // @[control.py:89:Tile.fir@577.4]
  wire [1:0] _T_618; // @[control.py:89:Tile.fir@578.4]
  wire  _T_636; // @[control.py:89:Tile.fir@596.4]
  wire  _T_637; // @[control.py:89:Tile.fir@597.4]
  wire  _T_638; // @[control.py:89:Tile.fir@598.4]
  wire  _T_639; // @[control.py:89:Tile.fir@599.4]
  wire  _T_640; // @[control.py:89:Tile.fir@600.4]
  wire  _T_641; // @[control.py:89:Tile.fir@601.4]
  wire  _T_642; // @[control.py:89:Tile.fir@602.4]
  wire  _T_643; // @[control.py:89:Tile.fir@603.4]
  wire  _T_644; // @[control.py:89:Tile.fir@604.4]
  wire  _T_645; // @[control.py:89:Tile.fir@605.4]
  wire  _T_646; // @[control.py:89:Tile.fir@606.4]
  wire  _T_647; // @[control.py:89:Tile.fir@607.4]
  wire  _T_648; // @[control.py:89:Tile.fir@608.4]
  wire  _T_649; // @[control.py:89:Tile.fir@609.4]
  wire  _T_650; // @[control.py:89:Tile.fir@610.4]
  wire  _T_651; // @[control.py:89:Tile.fir@611.4]
  wire  _T_652; // @[control.py:89:Tile.fir@612.4]
  wire  _T_653; // @[control.py:89:Tile.fir@613.4]
  wire  _T_654; // @[control.py:89:Tile.fir@614.4]
  wire  _T_655; // @[control.py:89:Tile.fir@615.4]
  wire  _T_656; // @[control.py:89:Tile.fir@616.4]
  wire [2:0] _T_659; // @[control.py:89:Tile.fir@619.4]
  wire [2:0] _T_660; // @[control.py:89:Tile.fir@620.4]
  wire [2:0] _T_661; // @[control.py:89:Tile.fir@621.4]
  wire [2:0] _T_662; // @[control.py:89:Tile.fir@622.4]
  wire [2:0] _T_663; // @[control.py:89:Tile.fir@623.4]
  wire [2:0] _T_664; // @[control.py:89:Tile.fir@624.4]
  wire [2:0] _T_665; // @[control.py:89:Tile.fir@625.4]
  wire [2:0] _T_666; // @[control.py:89:Tile.fir@626.4]
  wire [2:0] _T_667; // @[control.py:89:Tile.fir@627.4]
  wire [2:0] _T_668; // @[control.py:89:Tile.fir@628.4]
  wire [2:0] _T_669; // @[control.py:89:Tile.fir@629.4]
  wire [2:0] _T_670; // @[control.py:89:Tile.fir@630.4]
  wire [2:0] _T_671; // @[control.py:89:Tile.fir@631.4]
  wire [2:0] _T_672; // @[control.py:89:Tile.fir@632.4]
  wire [2:0] _T_673; // @[control.py:89:Tile.fir@633.4]
  wire [2:0] _T_674; // @[control.py:89:Tile.fir@634.4]
  wire [2:0] _T_675; // @[control.py:89:Tile.fir@635.4]
  wire [2:0] _T_676; // @[control.py:89:Tile.fir@636.4]
  wire [2:0] _T_677; // @[control.py:89:Tile.fir@637.4]
  wire [2:0] _T_678; // @[control.py:89:Tile.fir@638.4]
  wire [2:0] _T_679; // @[control.py:89:Tile.fir@639.4]
  wire [2:0] _T_680; // @[control.py:89:Tile.fir@640.4]
  wire [2:0] _T_681; // @[control.py:89:Tile.fir@641.4]
  wire [2:0] _T_682; // @[control.py:89:Tile.fir@642.4]
  wire [2:0] _T_683; // @[control.py:89:Tile.fir@643.4]
  wire [2:0] _T_684; // @[control.py:89:Tile.fir@644.4]
  wire [2:0] _T_685; // @[control.py:89:Tile.fir@645.4]
  wire [2:0] _T_686; // @[control.py:89:Tile.fir@646.4]
  wire [2:0] _T_687; // @[control.py:89:Tile.fir@647.4]
  wire [2:0] _T_688; // @[control.py:89:Tile.fir@648.4]
  wire [2:0] _T_689; // @[control.py:89:Tile.fir@649.4]
  wire [2:0] _T_690; // @[control.py:89:Tile.fir@650.4]
  wire [2:0] _T_691; // @[control.py:89:Tile.fir@651.4]
  wire [2:0] _T_692; // @[control.py:89:Tile.fir@652.4]
  wire [2:0] _T_693; // @[control.py:89:Tile.fir@653.4]
  wire [2:0] _T_694; // @[control.py:89:Tile.fir@654.4]
  wire  _T_701; // @[control.py:89:Tile.fir@661.4]
  wire  _T_702; // @[control.py:89:Tile.fir@662.4]
  wire  _T_703; // @[control.py:89:Tile.fir@663.4]
  wire  _T_704; // @[control.py:89:Tile.fir@664.4]
  wire  _T_705; // @[control.py:89:Tile.fir@665.4]
  wire  _T_706; // @[control.py:89:Tile.fir@666.4]
  wire  _T_707; // @[control.py:89:Tile.fir@667.4]
  wire  _T_708; // @[control.py:89:Tile.fir@668.4]
  wire  _T_709; // @[control.py:89:Tile.fir@669.4]
  wire  _T_710; // @[control.py:89:Tile.fir@670.4]
  wire  _T_711; // @[control.py:89:Tile.fir@671.4]
  wire  _T_712; // @[control.py:89:Tile.fir@672.4]
  wire  _T_713; // @[control.py:89:Tile.fir@673.4]
  wire  _T_714; // @[control.py:89:Tile.fir@674.4]
  wire  _T_715; // @[control.py:89:Tile.fir@675.4]
  wire  _T_716; // @[control.py:89:Tile.fir@676.4]
  wire  _T_717; // @[control.py:89:Tile.fir@677.4]
  wire  _T_718; // @[control.py:89:Tile.fir@678.4]
  wire  _T_719; // @[control.py:89:Tile.fir@679.4]
  wire  _T_720; // @[control.py:89:Tile.fir@680.4]
  wire  _T_721; // @[control.py:89:Tile.fir@681.4]
  wire  _T_722; // @[control.py:89:Tile.fir@682.4]
  wire  _T_723; // @[control.py:89:Tile.fir@683.4]
  wire  _T_724; // @[control.py:89:Tile.fir@684.4]
  wire  _T_725; // @[control.py:89:Tile.fir@685.4]
  wire  _T_726; // @[control.py:89:Tile.fir@686.4]
  wire  _T_727; // @[control.py:89:Tile.fir@687.4]
  wire  _T_728; // @[control.py:89:Tile.fir@688.4]
  wire  _T_729; // @[control.py:89:Tile.fir@689.4]
  wire  _T_730; // @[control.py:89:Tile.fir@690.4]
  wire  _T_731; // @[control.py:89:Tile.fir@691.4]
  wire  _T_732; // @[control.py:89:Tile.fir@692.4]
  assign _T_202 = io_inst & 32'hfe00707f; // @[listlookup.py:52:Tile.fir@162.4]
  assign _T_203 = _T_202 == 32'h33; // @[listlookup.py:52:Tile.fir@163.4]
  assign _T_205 = _T_202 == 32'h40000033; // @[listlookup.py:52:Tile.fir@165.4]
  assign _T_207 = _T_202 == 32'h7033; // @[listlookup.py:52:Tile.fir@167.4]
  assign _T_209 = _T_202 == 32'h6033; // @[listlookup.py:52:Tile.fir@169.4]
  assign _T_211 = _T_202 == 32'h4033; // @[listlookup.py:52:Tile.fir@171.4]
  assign _T_212 = io_inst & 32'h707f; // @[listlookup.py:52:Tile.fir@172.4]
  assign _T_213 = _T_212 == 32'h13; // @[listlookup.py:52:Tile.fir@173.4]
  assign _T_215 = _T_212 == 32'h7013; // @[listlookup.py:52:Tile.fir@175.4]
  assign _T_217 = _T_212 == 32'h6013; // @[listlookup.py:52:Tile.fir@177.4]
  assign _T_219 = _T_212 == 32'h4013; // @[listlookup.py:52:Tile.fir@179.4]
  assign _T_221 = _T_202 == 32'h1033; // @[listlookup.py:52:Tile.fir@181.4]
  assign _T_223 = _T_202 == 32'h5033; // @[listlookup.py:52:Tile.fir@183.4]
  assign _T_225 = _T_202 == 32'h40005033; // @[listlookup.py:52:Tile.fir@185.4]
  assign _T_227 = _T_202 == 32'h1013; // @[listlookup.py:52:Tile.fir@187.4]
  assign _T_229 = _T_202 == 32'h5013; // @[listlookup.py:52:Tile.fir@189.4]
  assign _T_231 = _T_202 == 32'h40005013; // @[listlookup.py:52:Tile.fir@191.4]
  assign _T_233 = _T_202 == 32'h2033; // @[listlookup.py:52:Tile.fir@193.4]
  assign _T_235 = _T_202 == 32'h3033; // @[listlookup.py:52:Tile.fir@195.4]
  assign _T_237 = _T_212 == 32'h2013; // @[listlookup.py:52:Tile.fir@197.4]
  assign _T_239 = _T_212 == 32'h3013; // @[listlookup.py:52:Tile.fir@199.4]
  assign _T_241 = _T_212 == 32'h2003; // @[listlookup.py:52:Tile.fir@201.4]
  assign _T_243 = _T_212 == 32'h1003; // @[listlookup.py:52:Tile.fir@203.4]
  assign _T_245 = _T_212 == 32'h3; // @[listlookup.py:52:Tile.fir@205.4]
  assign _T_247 = _T_212 == 32'h5003; // @[listlookup.py:52:Tile.fir@207.4]
  assign _T_249 = _T_212 == 32'h4003; // @[listlookup.py:52:Tile.fir@209.4]
  assign _T_251 = _T_212 == 32'h2023; // @[listlookup.py:52:Tile.fir@211.4]
  assign _T_253 = _T_212 == 32'h1023; // @[listlookup.py:52:Tile.fir@213.4]
  assign _T_255 = _T_212 == 32'h23; // @[listlookup.py:52:Tile.fir@215.4]
  assign _T_257 = _T_212 == 32'h63; // @[listlookup.py:52:Tile.fir@217.4]
  assign _T_259 = _T_212 == 32'h1063; // @[listlookup.py:52:Tile.fir@219.4]
  assign _T_261 = _T_212 == 32'h4063; // @[listlookup.py:52:Tile.fir@221.4]
  assign _T_263 = _T_212 == 32'h5063; // @[listlookup.py:52:Tile.fir@223.4]
  assign _T_265 = _T_212 == 32'h6063; // @[listlookup.py:52:Tile.fir@225.4]
  assign _T_267 = _T_212 == 32'h7063; // @[listlookup.py:52:Tile.fir@227.4]
  assign _T_268 = io_inst & 32'h7f; // @[listlookup.py:52:Tile.fir@228.4]
  assign _T_269 = _T_268 == 32'h6f; // @[listlookup.py:52:Tile.fir@229.4]
  assign _T_271 = _T_212 == 32'h67; // @[listlookup.py:52:Tile.fir@231.4]
  assign _T_273 = _T_268 == 32'h37; // @[listlookup.py:52:Tile.fir@233.4]
  assign _T_275 = _T_268 == 32'h17; // @[listlookup.py:52:Tile.fir@235.4]
  assign _T_280 = _T_273 ? 1'h1 : _T_275; // @[control.py:89:Tile.fir@240.4]
  assign _T_281 = _T_271 ? 1'h1 : _T_280; // @[control.py:89:Tile.fir@241.4]
  assign _T_282 = _T_269 ? 1'h1 : _T_281; // @[control.py:89:Tile.fir@242.4]
  assign _T_283 = _T_267 ? 1'h0 : _T_282; // @[control.py:89:Tile.fir@243.4]
  assign _T_284 = _T_265 ? 1'h0 : _T_283; // @[control.py:89:Tile.fir@244.4]
  assign _T_285 = _T_263 ? 1'h0 : _T_284; // @[control.py:89:Tile.fir@245.4]
  assign _T_286 = _T_261 ? 1'h0 : _T_285; // @[control.py:89:Tile.fir@246.4]
  assign _T_287 = _T_259 ? 1'h0 : _T_286; // @[control.py:89:Tile.fir@247.4]
  assign _T_288 = _T_257 ? 1'h0 : _T_287; // @[control.py:89:Tile.fir@248.4]
  assign _T_289 = _T_255 ? 1'h0 : _T_288; // @[control.py:89:Tile.fir@249.4]
  assign _T_290 = _T_253 ? 1'h0 : _T_289; // @[control.py:89:Tile.fir@250.4]
  assign _T_291 = _T_251 ? 1'h0 : _T_290; // @[control.py:89:Tile.fir@251.4]
  assign _T_292 = _T_249 ? 1'h1 : _T_291; // @[control.py:89:Tile.fir@252.4]
  assign _T_293 = _T_247 ? 1'h1 : _T_292; // @[control.py:89:Tile.fir@253.4]
  assign _T_294 = _T_245 ? 1'h1 : _T_293; // @[control.py:89:Tile.fir@254.4]
  assign _T_295 = _T_243 ? 1'h1 : _T_294; // @[control.py:89:Tile.fir@255.4]
  assign _T_296 = _T_241 ? 1'h1 : _T_295; // @[control.py:89:Tile.fir@256.4]
  assign _T_297 = _T_239 ? 1'h1 : _T_296; // @[control.py:89:Tile.fir@257.4]
  assign _T_298 = _T_237 ? 1'h1 : _T_297; // @[control.py:89:Tile.fir@258.4]
  assign _T_299 = _T_235 ? 1'h1 : _T_298; // @[control.py:89:Tile.fir@259.4]
  assign _T_300 = _T_233 ? 1'h1 : _T_299; // @[control.py:89:Tile.fir@260.4]
  assign _T_301 = _T_231 ? 1'h1 : _T_300; // @[control.py:89:Tile.fir@261.4]
  assign _T_302 = _T_229 ? 1'h1 : _T_301; // @[control.py:89:Tile.fir@262.4]
  assign _T_303 = _T_227 ? 1'h1 : _T_302; // @[control.py:89:Tile.fir@263.4]
  assign _T_304 = _T_225 ? 1'h1 : _T_303; // @[control.py:89:Tile.fir@264.4]
  assign _T_305 = _T_223 ? 1'h1 : _T_304; // @[control.py:89:Tile.fir@265.4]
  assign _T_306 = _T_221 ? 1'h1 : _T_305; // @[control.py:89:Tile.fir@266.4]
  assign _T_307 = _T_219 ? 1'h1 : _T_306; // @[control.py:89:Tile.fir@267.4]
  assign _T_308 = _T_217 ? 1'h1 : _T_307; // @[control.py:89:Tile.fir@268.4]
  assign _T_309 = _T_215 ? 1'h1 : _T_308; // @[control.py:89:Tile.fir@269.4]
  assign _T_310 = _T_213 ? 1'h1 : _T_309; // @[control.py:89:Tile.fir@270.4]
  assign _T_311 = _T_211 ? 1'h1 : _T_310; // @[control.py:89:Tile.fir@271.4]
  assign _T_312 = _T_209 ? 1'h1 : _T_311; // @[control.py:89:Tile.fir@272.4]
  assign _T_313 = _T_207 ? 1'h1 : _T_312; // @[control.py:89:Tile.fir@273.4]
  assign _T_314 = _T_205 ? 1'h1 : _T_313; // @[control.py:89:Tile.fir@274.4]
  assign _T_317 = _T_275 ? 3'h5 : 3'h0; // @[control.py:89:Tile.fir@277.4]
  assign _T_318 = _T_273 ? 3'h5 : _T_317; // @[control.py:89:Tile.fir@278.4]
  assign _T_319 = _T_271 ? 3'h2 : _T_318; // @[control.py:89:Tile.fir@279.4]
  assign _T_320 = _T_269 ? 3'h6 : _T_319; // @[control.py:89:Tile.fir@280.4]
  assign _T_321 = _T_267 ? 3'h4 : _T_320; // @[control.py:89:Tile.fir@281.4]
  assign _T_322 = _T_265 ? 3'h4 : _T_321; // @[control.py:89:Tile.fir@282.4]
  assign _T_323 = _T_263 ? 3'h4 : _T_322; // @[control.py:89:Tile.fir@283.4]
  assign _T_324 = _T_261 ? 3'h4 : _T_323; // @[control.py:89:Tile.fir@284.4]
  assign _T_325 = _T_259 ? 3'h4 : _T_324; // @[control.py:89:Tile.fir@285.4]
  assign _T_326 = _T_257 ? 3'h4 : _T_325; // @[control.py:89:Tile.fir@286.4]
  assign _T_327 = _T_255 ? 3'h3 : _T_326; // @[control.py:89:Tile.fir@287.4]
  assign _T_328 = _T_253 ? 3'h3 : _T_327; // @[control.py:89:Tile.fir@288.4]
  assign _T_329 = _T_251 ? 3'h3 : _T_328; // @[control.py:89:Tile.fir@289.4]
  assign _T_330 = _T_249 ? 3'h2 : _T_329; // @[control.py:89:Tile.fir@290.4]
  assign _T_331 = _T_247 ? 3'h2 : _T_330; // @[control.py:89:Tile.fir@291.4]
  assign _T_332 = _T_245 ? 3'h2 : _T_331; // @[control.py:89:Tile.fir@292.4]
  assign _T_333 = _T_243 ? 3'h2 : _T_332; // @[control.py:89:Tile.fir@293.4]
  assign _T_334 = _T_241 ? 3'h2 : _T_333; // @[control.py:89:Tile.fir@294.4]
  assign _T_335 = _T_239 ? 3'h2 : _T_334; // @[control.py:89:Tile.fir@295.4]
  assign _T_336 = _T_237 ? 3'h2 : _T_335; // @[control.py:89:Tile.fir@296.4]
  assign _T_337 = _T_235 ? 3'h1 : _T_336; // @[control.py:89:Tile.fir@297.4]
  assign _T_338 = _T_233 ? 3'h1 : _T_337; // @[control.py:89:Tile.fir@298.4]
  assign _T_339 = _T_231 ? 3'h2 : _T_338; // @[control.py:89:Tile.fir@299.4]
  assign _T_340 = _T_229 ? 3'h2 : _T_339; // @[control.py:89:Tile.fir@300.4]
  assign _T_341 = _T_227 ? 3'h2 : _T_340; // @[control.py:89:Tile.fir@301.4]
  assign _T_342 = _T_225 ? 3'h1 : _T_341; // @[control.py:89:Tile.fir@302.4]
  assign _T_343 = _T_223 ? 3'h1 : _T_342; // @[control.py:89:Tile.fir@303.4]
  assign _T_344 = _T_221 ? 3'h1 : _T_343; // @[control.py:89:Tile.fir@304.4]
  assign _T_345 = _T_219 ? 3'h2 : _T_344; // @[control.py:89:Tile.fir@305.4]
  assign _T_346 = _T_217 ? 3'h2 : _T_345; // @[control.py:89:Tile.fir@306.4]
  assign _T_347 = _T_215 ? 3'h2 : _T_346; // @[control.py:89:Tile.fir@307.4]
  assign _T_348 = _T_213 ? 3'h2 : _T_347; // @[control.py:89:Tile.fir@308.4]
  assign _T_349 = _T_211 ? 3'h1 : _T_348; // @[control.py:89:Tile.fir@309.4]
  assign _T_350 = _T_209 ? 3'h1 : _T_349; // @[control.py:89:Tile.fir@310.4]
  assign _T_351 = _T_207 ? 3'h1 : _T_350; // @[control.py:89:Tile.fir@311.4]
  assign _T_352 = _T_205 ? 3'h1 : _T_351; // @[control.py:89:Tile.fir@312.4]
  assign _T_366 = _T_253 ? 1'h1 : _T_255; // @[control.py:89:Tile.fir@326.4]
  assign _T_367 = _T_251 ? 1'h1 : _T_366; // @[control.py:89:Tile.fir@327.4]
  assign _T_368 = _T_249 ? 1'h1 : _T_367; // @[control.py:89:Tile.fir@328.4]
  assign _T_369 = _T_247 ? 1'h1 : _T_368; // @[control.py:89:Tile.fir@329.4]
  assign _T_370 = _T_245 ? 1'h1 : _T_369; // @[control.py:89:Tile.fir@330.4]
  assign _T_371 = _T_243 ? 1'h1 : _T_370; // @[control.py:89:Tile.fir@331.4]
  assign _T_372 = _T_241 ? 1'h1 : _T_371; // @[control.py:89:Tile.fir@332.4]
  assign _T_373 = _T_239 ? 1'h1 : _T_372; // @[control.py:89:Tile.fir@333.4]
  assign _T_374 = _T_237 ? 1'h1 : _T_373; // @[control.py:89:Tile.fir@334.4]
  assign _T_375 = _T_235 ? 1'h0 : _T_374; // @[control.py:89:Tile.fir@335.4]
  assign _T_376 = _T_233 ? 1'h0 : _T_375; // @[control.py:89:Tile.fir@336.4]
  assign _T_377 = _T_231 ? 1'h1 : _T_376; // @[control.py:89:Tile.fir@337.4]
  assign _T_378 = _T_229 ? 1'h1 : _T_377; // @[control.py:89:Tile.fir@338.4]
  assign _T_379 = _T_227 ? 1'h1 : _T_378; // @[control.py:89:Tile.fir@339.4]
  assign _T_380 = _T_225 ? 1'h0 : _T_379; // @[control.py:89:Tile.fir@340.4]
  assign _T_381 = _T_223 ? 1'h0 : _T_380; // @[control.py:89:Tile.fir@341.4]
  assign _T_382 = _T_221 ? 1'h0 : _T_381; // @[control.py:89:Tile.fir@342.4]
  assign _T_383 = _T_219 ? 1'h1 : _T_382; // @[control.py:89:Tile.fir@343.4]
  assign _T_384 = _T_217 ? 1'h1 : _T_383; // @[control.py:89:Tile.fir@344.4]
  assign _T_385 = _T_215 ? 1'h1 : _T_384; // @[control.py:89:Tile.fir@345.4]
  assign _T_386 = _T_213 ? 1'h1 : _T_385; // @[control.py:89:Tile.fir@346.4]
  assign _T_387 = _T_211 ? 1'h0 : _T_386; // @[control.py:89:Tile.fir@347.4]
  assign _T_388 = _T_209 ? 1'h0 : _T_387; // @[control.py:89:Tile.fir@348.4]
  assign _T_389 = _T_207 ? 1'h0 : _T_388; // @[control.py:89:Tile.fir@349.4]
  assign _T_390 = _T_205 ? 1'h0 : _T_389; // @[control.py:89:Tile.fir@350.4]
  assign _T_393 = _T_275 ? 5'h0 : 5'h10; // @[control.py:89:Tile.fir@353.4]
  assign _T_394 = _T_273 ? 5'h0 : _T_393; // @[control.py:89:Tile.fir@354.4]
  assign _T_395 = _T_271 ? 5'h0 : _T_394; // @[control.py:89:Tile.fir@355.4]
  assign _T_396 = _T_269 ? 5'h0 : _T_395; // @[control.py:89:Tile.fir@356.4]
  assign _T_397 = _T_267 ? 5'hf : _T_396; // @[control.py:89:Tile.fir@357.4]
  assign _T_398 = _T_265 ? 5'he : _T_397; // @[control.py:89:Tile.fir@358.4]
  assign _T_399 = _T_263 ? 5'hd : _T_398; // @[control.py:89:Tile.fir@359.4]
  assign _T_400 = _T_261 ? 5'hc : _T_399; // @[control.py:89:Tile.fir@360.4]
  assign _T_401 = _T_259 ? 5'hb : _T_400; // @[control.py:89:Tile.fir@361.4]
  assign _T_402 = _T_257 ? 5'ha : _T_401; // @[control.py:89:Tile.fir@362.4]
  assign _T_403 = _T_255 ? 5'h0 : _T_402; // @[control.py:89:Tile.fir@363.4]
  assign _T_404 = _T_253 ? 5'h0 : _T_403; // @[control.py:89:Tile.fir@364.4]
  assign _T_405 = _T_251 ? 5'h0 : _T_404; // @[control.py:89:Tile.fir@365.4]
  assign _T_406 = _T_249 ? 5'h0 : _T_405; // @[control.py:89:Tile.fir@366.4]
  assign _T_407 = _T_247 ? 5'h0 : _T_406; // @[control.py:89:Tile.fir@367.4]
  assign _T_408 = _T_245 ? 5'h0 : _T_407; // @[control.py:89:Tile.fir@368.4]
  assign _T_409 = _T_243 ? 5'h0 : _T_408; // @[control.py:89:Tile.fir@369.4]
  assign _T_410 = _T_241 ? 5'h0 : _T_409; // @[control.py:89:Tile.fir@370.4]
  assign _T_411 = _T_239 ? 5'h9 : _T_410; // @[control.py:89:Tile.fir@371.4]
  assign _T_412 = _T_237 ? 5'h8 : _T_411; // @[control.py:89:Tile.fir@372.4]
  assign _T_413 = _T_235 ? 5'h9 : _T_412; // @[control.py:89:Tile.fir@373.4]
  assign _T_414 = _T_233 ? 5'h8 : _T_413; // @[control.py:89:Tile.fir@374.4]
  assign _T_415 = _T_231 ? 5'h7 : _T_414; // @[control.py:89:Tile.fir@375.4]
  assign _T_416 = _T_229 ? 5'h6 : _T_415; // @[control.py:89:Tile.fir@376.4]
  assign _T_417 = _T_227 ? 5'h5 : _T_416; // @[control.py:89:Tile.fir@377.4]
  assign _T_418 = _T_225 ? 5'h7 : _T_417; // @[control.py:89:Tile.fir@378.4]
  assign _T_419 = _T_223 ? 5'h6 : _T_418; // @[control.py:89:Tile.fir@379.4]
  assign _T_420 = _T_221 ? 5'h5 : _T_419; // @[control.py:89:Tile.fir@380.4]
  assign _T_421 = _T_219 ? 5'h4 : _T_420; // @[control.py:89:Tile.fir@381.4]
  assign _T_422 = _T_217 ? 5'h3 : _T_421; // @[control.py:89:Tile.fir@382.4]
  assign _T_423 = _T_215 ? 5'h2 : _T_422; // @[control.py:89:Tile.fir@383.4]
  assign _T_424 = _T_213 ? 5'h0 : _T_423; // @[control.py:89:Tile.fir@384.4]
  assign _T_425 = _T_211 ? 5'h4 : _T_424; // @[control.py:89:Tile.fir@385.4]
  assign _T_426 = _T_209 ? 5'h3 : _T_425; // @[control.py:89:Tile.fir@386.4]
  assign _T_427 = _T_207 ? 5'h2 : _T_426; // @[control.py:89:Tile.fir@387.4]
  assign _T_428 = _T_205 ? 5'h1 : _T_427; // @[control.py:89:Tile.fir@388.4]
  assign _T_434 = _T_269 ? 1'h1 : _T_271; // @[control.py:89:Tile.fir@394.4]
  assign _T_435 = _T_267 ? 1'h1 : _T_434; // @[control.py:89:Tile.fir@395.4]
  assign _T_436 = _T_265 ? 1'h1 : _T_435; // @[control.py:89:Tile.fir@396.4]
  assign _T_437 = _T_263 ? 1'h1 : _T_436; // @[control.py:89:Tile.fir@397.4]
  assign _T_438 = _T_261 ? 1'h1 : _T_437; // @[control.py:89:Tile.fir@398.4]
  assign _T_439 = _T_259 ? 1'h1 : _T_438; // @[control.py:89:Tile.fir@399.4]
  assign _T_440 = _T_257 ? 1'h1 : _T_439; // @[control.py:89:Tile.fir@400.4]
  assign _T_441 = _T_255 ? 1'h0 : _T_440; // @[control.py:89:Tile.fir@401.4]
  assign _T_442 = _T_253 ? 1'h0 : _T_441; // @[control.py:89:Tile.fir@402.4]
  assign _T_443 = _T_251 ? 1'h0 : _T_442; // @[control.py:89:Tile.fir@403.4]
  assign _T_444 = _T_249 ? 1'h0 : _T_443; // @[control.py:89:Tile.fir@404.4]
  assign _T_445 = _T_247 ? 1'h0 : _T_444; // @[control.py:89:Tile.fir@405.4]
  assign _T_446 = _T_245 ? 1'h0 : _T_445; // @[control.py:89:Tile.fir@406.4]
  assign _T_447 = _T_243 ? 1'h0 : _T_446; // @[control.py:89:Tile.fir@407.4]
  assign _T_448 = _T_241 ? 1'h0 : _T_447; // @[control.py:89:Tile.fir@408.4]
  assign _T_449 = _T_239 ? 1'h0 : _T_448; // @[control.py:89:Tile.fir@409.4]
  assign _T_450 = _T_237 ? 1'h0 : _T_449; // @[control.py:89:Tile.fir@410.4]
  assign _T_451 = _T_235 ? 1'h0 : _T_450; // @[control.py:89:Tile.fir@411.4]
  assign _T_452 = _T_233 ? 1'h0 : _T_451; // @[control.py:89:Tile.fir@412.4]
  assign _T_453 = _T_231 ? 1'h0 : _T_452; // @[control.py:89:Tile.fir@413.4]
  assign _T_454 = _T_229 ? 1'h0 : _T_453; // @[control.py:89:Tile.fir@414.4]
  assign _T_455 = _T_227 ? 1'h0 : _T_454; // @[control.py:89:Tile.fir@415.4]
  assign _T_456 = _T_225 ? 1'h0 : _T_455; // @[control.py:89:Tile.fir@416.4]
  assign _T_457 = _T_223 ? 1'h0 : _T_456; // @[control.py:89:Tile.fir@417.4]
  assign _T_458 = _T_221 ? 1'h0 : _T_457; // @[control.py:89:Tile.fir@418.4]
  assign _T_459 = _T_219 ? 1'h0 : _T_458; // @[control.py:89:Tile.fir@419.4]
  assign _T_460 = _T_217 ? 1'h0 : _T_459; // @[control.py:89:Tile.fir@420.4]
  assign _T_461 = _T_215 ? 1'h0 : _T_460; // @[control.py:89:Tile.fir@421.4]
  assign _T_462 = _T_213 ? 1'h0 : _T_461; // @[control.py:89:Tile.fir@422.4]
  assign _T_463 = _T_211 ? 1'h0 : _T_462; // @[control.py:89:Tile.fir@423.4]
  assign _T_464 = _T_209 ? 1'h0 : _T_463; // @[control.py:89:Tile.fir@424.4]
  assign _T_465 = _T_207 ? 1'h0 : _T_464; // @[control.py:89:Tile.fir@425.4]
  assign _T_466 = _T_205 ? 1'h0 : _T_465; // @[control.py:89:Tile.fir@426.4]
  assign _T_472 = _T_269 ? 1'h0 : _T_271; // @[control.py:89:Tile.fir@432.4]
  assign _T_473 = _T_267 ? 1'h0 : _T_472; // @[control.py:89:Tile.fir@433.4]
  assign _T_474 = _T_265 ? 1'h0 : _T_473; // @[control.py:89:Tile.fir@434.4]
  assign _T_475 = _T_263 ? 1'h0 : _T_474; // @[control.py:89:Tile.fir@435.4]
  assign _T_476 = _T_261 ? 1'h0 : _T_475; // @[control.py:89:Tile.fir@436.4]
  assign _T_477 = _T_259 ? 1'h0 : _T_476; // @[control.py:89:Tile.fir@437.4]
  assign _T_478 = _T_257 ? 1'h0 : _T_477; // @[control.py:89:Tile.fir@438.4]
  assign _T_479 = _T_255 ? 1'h0 : _T_478; // @[control.py:89:Tile.fir@439.4]
  assign _T_480 = _T_253 ? 1'h0 : _T_479; // @[control.py:89:Tile.fir@440.4]
  assign _T_481 = _T_251 ? 1'h0 : _T_480; // @[control.py:89:Tile.fir@441.4]
  assign _T_482 = _T_249 ? 1'h0 : _T_481; // @[control.py:89:Tile.fir@442.4]
  assign _T_483 = _T_247 ? 1'h0 : _T_482; // @[control.py:89:Tile.fir@443.4]
  assign _T_484 = _T_245 ? 1'h0 : _T_483; // @[control.py:89:Tile.fir@444.4]
  assign _T_485 = _T_243 ? 1'h0 : _T_484; // @[control.py:89:Tile.fir@445.4]
  assign _T_486 = _T_241 ? 1'h0 : _T_485; // @[control.py:89:Tile.fir@446.4]
  assign _T_487 = _T_239 ? 1'h0 : _T_486; // @[control.py:89:Tile.fir@447.4]
  assign _T_488 = _T_237 ? 1'h0 : _T_487; // @[control.py:89:Tile.fir@448.4]
  assign _T_489 = _T_235 ? 1'h0 : _T_488; // @[control.py:89:Tile.fir@449.4]
  assign _T_490 = _T_233 ? 1'h0 : _T_489; // @[control.py:89:Tile.fir@450.4]
  assign _T_491 = _T_231 ? 1'h0 : _T_490; // @[control.py:89:Tile.fir@451.4]
  assign _T_492 = _T_229 ? 1'h0 : _T_491; // @[control.py:89:Tile.fir@452.4]
  assign _T_493 = _T_227 ? 1'h0 : _T_492; // @[control.py:89:Tile.fir@453.4]
  assign _T_494 = _T_225 ? 1'h0 : _T_493; // @[control.py:89:Tile.fir@454.4]
  assign _T_495 = _T_223 ? 1'h0 : _T_494; // @[control.py:89:Tile.fir@455.4]
  assign _T_496 = _T_221 ? 1'h0 : _T_495; // @[control.py:89:Tile.fir@456.4]
  assign _T_497 = _T_219 ? 1'h0 : _T_496; // @[control.py:89:Tile.fir@457.4]
  assign _T_498 = _T_217 ? 1'h0 : _T_497; // @[control.py:89:Tile.fir@458.4]
  assign _T_499 = _T_215 ? 1'h0 : _T_498; // @[control.py:89:Tile.fir@459.4]
  assign _T_500 = _T_213 ? 1'h0 : _T_499; // @[control.py:89:Tile.fir@460.4]
  assign _T_501 = _T_211 ? 1'h0 : _T_500; // @[control.py:89:Tile.fir@461.4]
  assign _T_502 = _T_209 ? 1'h0 : _T_501; // @[control.py:89:Tile.fir@462.4]
  assign _T_503 = _T_207 ? 1'h0 : _T_502; // @[control.py:89:Tile.fir@463.4]
  assign _T_504 = _T_205 ? 1'h0 : _T_503; // @[control.py:89:Tile.fir@464.4]
  assign _T_521 = _T_247 ? 1'h1 : _T_249; // @[control.py:89:Tile.fir@481.4]
  assign _T_522 = _T_245 ? 1'h1 : _T_521; // @[control.py:89:Tile.fir@482.4]
  assign _T_523 = _T_243 ? 1'h1 : _T_522; // @[control.py:89:Tile.fir@483.4]
  assign _T_524 = _T_241 ? 1'h1 : _T_523; // @[control.py:89:Tile.fir@484.4]
  assign _T_525 = _T_239 ? 1'h0 : _T_524; // @[control.py:89:Tile.fir@485.4]
  assign _T_526 = _T_237 ? 1'h0 : _T_525; // @[control.py:89:Tile.fir@486.4]
  assign _T_527 = _T_235 ? 1'h0 : _T_526; // @[control.py:89:Tile.fir@487.4]
  assign _T_528 = _T_233 ? 1'h0 : _T_527; // @[control.py:89:Tile.fir@488.4]
  assign _T_529 = _T_231 ? 1'h0 : _T_528; // @[control.py:89:Tile.fir@489.4]
  assign _T_530 = _T_229 ? 1'h0 : _T_529; // @[control.py:89:Tile.fir@490.4]
  assign _T_531 = _T_227 ? 1'h0 : _T_530; // @[control.py:89:Tile.fir@491.4]
  assign _T_532 = _T_225 ? 1'h0 : _T_531; // @[control.py:89:Tile.fir@492.4]
  assign _T_533 = _T_223 ? 1'h0 : _T_532; // @[control.py:89:Tile.fir@493.4]
  assign _T_534 = _T_221 ? 1'h0 : _T_533; // @[control.py:89:Tile.fir@494.4]
  assign _T_535 = _T_219 ? 1'h0 : _T_534; // @[control.py:89:Tile.fir@495.4]
  assign _T_536 = _T_217 ? 1'h0 : _T_535; // @[control.py:89:Tile.fir@496.4]
  assign _T_537 = _T_215 ? 1'h0 : _T_536; // @[control.py:89:Tile.fir@497.4]
  assign _T_538 = _T_213 ? 1'h0 : _T_537; // @[control.py:89:Tile.fir@498.4]
  assign _T_539 = _T_211 ? 1'h0 : _T_538; // @[control.py:89:Tile.fir@499.4]
  assign _T_540 = _T_209 ? 1'h0 : _T_539; // @[control.py:89:Tile.fir@500.4]
  assign _T_541 = _T_207 ? 1'h0 : _T_540; // @[control.py:89:Tile.fir@501.4]
  assign _T_542 = _T_205 ? 1'h0 : _T_541; // @[control.py:89:Tile.fir@502.4]
  assign _T_558 = _T_249 ? 1'h0 : _T_367; // @[control.py:89:Tile.fir@518.4]
  assign _T_559 = _T_247 ? 1'h0 : _T_558; // @[control.py:89:Tile.fir@519.4]
  assign _T_560 = _T_245 ? 1'h0 : _T_559; // @[control.py:89:Tile.fir@520.4]
  assign _T_561 = _T_243 ? 1'h0 : _T_560; // @[control.py:89:Tile.fir@521.4]
  assign _T_562 = _T_241 ? 1'h0 : _T_561; // @[control.py:89:Tile.fir@522.4]
  assign _T_563 = _T_239 ? 1'h0 : _T_562; // @[control.py:89:Tile.fir@523.4]
  assign _T_564 = _T_237 ? 1'h0 : _T_563; // @[control.py:89:Tile.fir@524.4]
  assign _T_565 = _T_235 ? 1'h0 : _T_564; // @[control.py:89:Tile.fir@525.4]
  assign _T_566 = _T_233 ? 1'h0 : _T_565; // @[control.py:89:Tile.fir@526.4]
  assign _T_567 = _T_231 ? 1'h0 : _T_566; // @[control.py:89:Tile.fir@527.4]
  assign _T_568 = _T_229 ? 1'h0 : _T_567; // @[control.py:89:Tile.fir@528.4]
  assign _T_569 = _T_227 ? 1'h0 : _T_568; // @[control.py:89:Tile.fir@529.4]
  assign _T_570 = _T_225 ? 1'h0 : _T_569; // @[control.py:89:Tile.fir@530.4]
  assign _T_571 = _T_223 ? 1'h0 : _T_570; // @[control.py:89:Tile.fir@531.4]
  assign _T_572 = _T_221 ? 1'h0 : _T_571; // @[control.py:89:Tile.fir@532.4]
  assign _T_573 = _T_219 ? 1'h0 : _T_572; // @[control.py:89:Tile.fir@533.4]
  assign _T_574 = _T_217 ? 1'h0 : _T_573; // @[control.py:89:Tile.fir@534.4]
  assign _T_575 = _T_215 ? 1'h0 : _T_574; // @[control.py:89:Tile.fir@535.4]
  assign _T_576 = _T_213 ? 1'h0 : _T_575; // @[control.py:89:Tile.fir@536.4]
  assign _T_577 = _T_211 ? 1'h0 : _T_576; // @[control.py:89:Tile.fir@537.4]
  assign _T_578 = _T_209 ? 1'h0 : _T_577; // @[control.py:89:Tile.fir@538.4]
  assign _T_579 = _T_207 ? 1'h0 : _T_578; // @[control.py:89:Tile.fir@539.4]
  assign _T_580 = _T_205 ? 1'h0 : _T_579; // @[control.py:89:Tile.fir@540.4]
  assign _T_593 = _T_255 ? 2'h2 : 2'h0; // @[control.py:89:Tile.fir@553.4]
  assign _T_594 = _T_253 ? 2'h1 : _T_593; // @[control.py:89:Tile.fir@554.4]
  assign _T_595 = _T_251 ? 2'h0 : _T_594; // @[control.py:89:Tile.fir@555.4]
  assign _T_596 = _T_249 ? 2'h2 : _T_595; // @[control.py:89:Tile.fir@556.4]
  assign _T_597 = _T_247 ? 2'h1 : _T_596; // @[control.py:89:Tile.fir@557.4]
  assign _T_598 = _T_245 ? 2'h2 : _T_597; // @[control.py:89:Tile.fir@558.4]
  assign _T_599 = _T_243 ? 2'h1 : _T_598; // @[control.py:89:Tile.fir@559.4]
  assign _T_600 = _T_241 ? 2'h0 : _T_599; // @[control.py:89:Tile.fir@560.4]
  assign _T_601 = _T_239 ? 2'h0 : _T_600; // @[control.py:89:Tile.fir@561.4]
  assign _T_602 = _T_237 ? 2'h0 : _T_601; // @[control.py:89:Tile.fir@562.4]
  assign _T_603 = _T_235 ? 2'h0 : _T_602; // @[control.py:89:Tile.fir@563.4]
  assign _T_604 = _T_233 ? 2'h0 : _T_603; // @[control.py:89:Tile.fir@564.4]
  assign _T_605 = _T_231 ? 2'h0 : _T_604; // @[control.py:89:Tile.fir@565.4]
  assign _T_606 = _T_229 ? 2'h0 : _T_605; // @[control.py:89:Tile.fir@566.4]
  assign _T_607 = _T_227 ? 2'h0 : _T_606; // @[control.py:89:Tile.fir@567.4]
  assign _T_608 = _T_225 ? 2'h0 : _T_607; // @[control.py:89:Tile.fir@568.4]
  assign _T_609 = _T_223 ? 2'h0 : _T_608; // @[control.py:89:Tile.fir@569.4]
  assign _T_610 = _T_221 ? 2'h0 : _T_609; // @[control.py:89:Tile.fir@570.4]
  assign _T_611 = _T_219 ? 2'h0 : _T_610; // @[control.py:89:Tile.fir@571.4]
  assign _T_612 = _T_217 ? 2'h0 : _T_611; // @[control.py:89:Tile.fir@572.4]
  assign _T_613 = _T_215 ? 2'h0 : _T_612; // @[control.py:89:Tile.fir@573.4]
  assign _T_614 = _T_213 ? 2'h0 : _T_613; // @[control.py:89:Tile.fir@574.4]
  assign _T_615 = _T_211 ? 2'h0 : _T_614; // @[control.py:89:Tile.fir@575.4]
  assign _T_616 = _T_209 ? 2'h0 : _T_615; // @[control.py:89:Tile.fir@576.4]
  assign _T_617 = _T_207 ? 2'h0 : _T_616; // @[control.py:89:Tile.fir@577.4]
  assign _T_618 = _T_205 ? 2'h0 : _T_617; // @[control.py:89:Tile.fir@578.4]
  assign _T_636 = _T_245 ? 1'h0 : _T_521; // @[control.py:89:Tile.fir@596.4]
  assign _T_637 = _T_243 ? 1'h0 : _T_636; // @[control.py:89:Tile.fir@597.4]
  assign _T_638 = _T_241 ? 1'h0 : _T_637; // @[control.py:89:Tile.fir@598.4]
  assign _T_639 = _T_239 ? 1'h0 : _T_638; // @[control.py:89:Tile.fir@599.4]
  assign _T_640 = _T_237 ? 1'h0 : _T_639; // @[control.py:89:Tile.fir@600.4]
  assign _T_641 = _T_235 ? 1'h0 : _T_640; // @[control.py:89:Tile.fir@601.4]
  assign _T_642 = _T_233 ? 1'h0 : _T_641; // @[control.py:89:Tile.fir@602.4]
  assign _T_643 = _T_231 ? 1'h0 : _T_642; // @[control.py:89:Tile.fir@603.4]
  assign _T_644 = _T_229 ? 1'h0 : _T_643; // @[control.py:89:Tile.fir@604.4]
  assign _T_645 = _T_227 ? 1'h0 : _T_644; // @[control.py:89:Tile.fir@605.4]
  assign _T_646 = _T_225 ? 1'h0 : _T_645; // @[control.py:89:Tile.fir@606.4]
  assign _T_647 = _T_223 ? 1'h0 : _T_646; // @[control.py:89:Tile.fir@607.4]
  assign _T_648 = _T_221 ? 1'h0 : _T_647; // @[control.py:89:Tile.fir@608.4]
  assign _T_649 = _T_219 ? 1'h0 : _T_648; // @[control.py:89:Tile.fir@609.4]
  assign _T_650 = _T_217 ? 1'h0 : _T_649; // @[control.py:89:Tile.fir@610.4]
  assign _T_651 = _T_215 ? 1'h0 : _T_650; // @[control.py:89:Tile.fir@611.4]
  assign _T_652 = _T_213 ? 1'h0 : _T_651; // @[control.py:89:Tile.fir@612.4]
  assign _T_653 = _T_211 ? 1'h0 : _T_652; // @[control.py:89:Tile.fir@613.4]
  assign _T_654 = _T_209 ? 1'h0 : _T_653; // @[control.py:89:Tile.fir@614.4]
  assign _T_655 = _T_207 ? 1'h0 : _T_654; // @[control.py:89:Tile.fir@615.4]
  assign _T_656 = _T_205 ? 1'h0 : _T_655; // @[control.py:89:Tile.fir@616.4]
  assign _T_659 = _T_275 ? 3'h4 : 3'h0; // @[control.py:89:Tile.fir@619.4]
  assign _T_660 = _T_273 ? 3'h3 : _T_659; // @[control.py:89:Tile.fir@620.4]
  assign _T_661 = _T_271 ? 3'h2 : _T_660; // @[control.py:89:Tile.fir@621.4]
  assign _T_662 = _T_269 ? 3'h2 : _T_661; // @[control.py:89:Tile.fir@622.4]
  assign _T_663 = _T_267 ? 3'h0 : _T_662; // @[control.py:89:Tile.fir@623.4]
  assign _T_664 = _T_265 ? 3'h0 : _T_663; // @[control.py:89:Tile.fir@624.4]
  assign _T_665 = _T_263 ? 3'h0 : _T_664; // @[control.py:89:Tile.fir@625.4]
  assign _T_666 = _T_261 ? 3'h0 : _T_665; // @[control.py:89:Tile.fir@626.4]
  assign _T_667 = _T_259 ? 3'h0 : _T_666; // @[control.py:89:Tile.fir@627.4]
  assign _T_668 = _T_257 ? 3'h0 : _T_667; // @[control.py:89:Tile.fir@628.4]
  assign _T_669 = _T_255 ? 3'h0 : _T_668; // @[control.py:89:Tile.fir@629.4]
  assign _T_670 = _T_253 ? 3'h0 : _T_669; // @[control.py:89:Tile.fir@630.4]
  assign _T_671 = _T_251 ? 3'h0 : _T_670; // @[control.py:89:Tile.fir@631.4]
  assign _T_672 = _T_249 ? 3'h1 : _T_671; // @[control.py:89:Tile.fir@632.4]
  assign _T_673 = _T_247 ? 3'h1 : _T_672; // @[control.py:89:Tile.fir@633.4]
  assign _T_674 = _T_245 ? 3'h1 : _T_673; // @[control.py:89:Tile.fir@634.4]
  assign _T_675 = _T_243 ? 3'h1 : _T_674; // @[control.py:89:Tile.fir@635.4]
  assign _T_676 = _T_241 ? 3'h1 : _T_675; // @[control.py:89:Tile.fir@636.4]
  assign _T_677 = _T_239 ? 3'h0 : _T_676; // @[control.py:89:Tile.fir@637.4]
  assign _T_678 = _T_237 ? 3'h0 : _T_677; // @[control.py:89:Tile.fir@638.4]
  assign _T_679 = _T_235 ? 3'h0 : _T_678; // @[control.py:89:Tile.fir@639.4]
  assign _T_680 = _T_233 ? 3'h0 : _T_679; // @[control.py:89:Tile.fir@640.4]
  assign _T_681 = _T_231 ? 3'h0 : _T_680; // @[control.py:89:Tile.fir@641.4]
  assign _T_682 = _T_229 ? 3'h0 : _T_681; // @[control.py:89:Tile.fir@642.4]
  assign _T_683 = _T_227 ? 3'h0 : _T_682; // @[control.py:89:Tile.fir@643.4]
  assign _T_684 = _T_225 ? 3'h0 : _T_683; // @[control.py:89:Tile.fir@644.4]
  assign _T_685 = _T_223 ? 3'h0 : _T_684; // @[control.py:89:Tile.fir@645.4]
  assign _T_686 = _T_221 ? 3'h0 : _T_685; // @[control.py:89:Tile.fir@646.4]
  assign _T_687 = _T_219 ? 3'h0 : _T_686; // @[control.py:89:Tile.fir@647.4]
  assign _T_688 = _T_217 ? 3'h0 : _T_687; // @[control.py:89:Tile.fir@648.4]
  assign _T_689 = _T_215 ? 3'h0 : _T_688; // @[control.py:89:Tile.fir@649.4]
  assign _T_690 = _T_213 ? 3'h0 : _T_689; // @[control.py:89:Tile.fir@650.4]
  assign _T_691 = _T_211 ? 3'h0 : _T_690; // @[control.py:89:Tile.fir@651.4]
  assign _T_692 = _T_209 ? 3'h0 : _T_691; // @[control.py:89:Tile.fir@652.4]
  assign _T_693 = _T_207 ? 3'h0 : _T_692; // @[control.py:89:Tile.fir@653.4]
  assign _T_694 = _T_205 ? 3'h0 : _T_693; // @[control.py:89:Tile.fir@654.4]
  assign _T_701 = _T_267 ? 1'h0 : _T_434; // @[control.py:89:Tile.fir@661.4]
  assign _T_702 = _T_265 ? 1'h0 : _T_701; // @[control.py:89:Tile.fir@662.4]
  assign _T_703 = _T_263 ? 1'h0 : _T_702; // @[control.py:89:Tile.fir@663.4]
  assign _T_704 = _T_261 ? 1'h0 : _T_703; // @[control.py:89:Tile.fir@664.4]
  assign _T_705 = _T_259 ? 1'h0 : _T_704; // @[control.py:89:Tile.fir@665.4]
  assign _T_706 = _T_257 ? 1'h0 : _T_705; // @[control.py:89:Tile.fir@666.4]
  assign _T_707 = _T_255 ? 1'h0 : _T_706; // @[control.py:89:Tile.fir@667.4]
  assign _T_708 = _T_253 ? 1'h0 : _T_707; // @[control.py:89:Tile.fir@668.4]
  assign _T_709 = _T_251 ? 1'h0 : _T_708; // @[control.py:89:Tile.fir@669.4]
  assign _T_710 = _T_249 ? 1'h0 : _T_709; // @[control.py:89:Tile.fir@670.4]
  assign _T_711 = _T_247 ? 1'h0 : _T_710; // @[control.py:89:Tile.fir@671.4]
  assign _T_712 = _T_245 ? 1'h0 : _T_711; // @[control.py:89:Tile.fir@672.4]
  assign _T_713 = _T_243 ? 1'h0 : _T_712; // @[control.py:89:Tile.fir@673.4]
  assign _T_714 = _T_241 ? 1'h0 : _T_713; // @[control.py:89:Tile.fir@674.4]
  assign _T_715 = _T_239 ? 1'h0 : _T_714; // @[control.py:89:Tile.fir@675.4]
  assign _T_716 = _T_237 ? 1'h0 : _T_715; // @[control.py:89:Tile.fir@676.4]
  assign _T_717 = _T_235 ? 1'h0 : _T_716; // @[control.py:89:Tile.fir@677.4]
  assign _T_718 = _T_233 ? 1'h0 : _T_717; // @[control.py:89:Tile.fir@678.4]
  assign _T_719 = _T_231 ? 1'h0 : _T_718; // @[control.py:89:Tile.fir@679.4]
  assign _T_720 = _T_229 ? 1'h0 : _T_719; // @[control.py:89:Tile.fir@680.4]
  assign _T_721 = _T_227 ? 1'h0 : _T_720; // @[control.py:89:Tile.fir@681.4]
  assign _T_722 = _T_225 ? 1'h0 : _T_721; // @[control.py:89:Tile.fir@682.4]
  assign _T_723 = _T_223 ? 1'h0 : _T_722; // @[control.py:89:Tile.fir@683.4]
  assign _T_724 = _T_221 ? 1'h0 : _T_723; // @[control.py:89:Tile.fir@684.4]
  assign _T_725 = _T_219 ? 1'h0 : _T_724; // @[control.py:89:Tile.fir@685.4]
  assign _T_726 = _T_217 ? 1'h0 : _T_725; // @[control.py:89:Tile.fir@686.4]
  assign _T_727 = _T_215 ? 1'h0 : _T_726; // @[control.py:89:Tile.fir@687.4]
  assign _T_728 = _T_213 ? 1'h0 : _T_727; // @[control.py:89:Tile.fir@688.4]
  assign _T_729 = _T_211 ? 1'h0 : _T_728; // @[control.py:89:Tile.fir@689.4]
  assign _T_730 = _T_209 ? 1'h0 : _T_729; // @[control.py:89:Tile.fir@690.4]
  assign _T_731 = _T_207 ? 1'h0 : _T_730; // @[control.py:89:Tile.fir@691.4]
  assign _T_732 = _T_205 ? 1'h0 : _T_731; // @[control.py:89:Tile.fir@692.4]
  assign io_Reg_Write = _T_203 ? 1'h1 : _T_314; // @[control.py:108:Tile.fir@704.4]
  assign io_Imm_Sel = _T_203 ? 3'h1 : _T_352; // @[control.py:92:Tile.fir@694.4]
  assign io_ALU_Src = _T_203 ? 1'h0 : _T_390; // @[control.py:95:Tile.fir@695.4]
  assign io_ALUOp = _T_203 ? 5'h0 : _T_428; // @[control.py:96:Tile.fir@696.4]
  assign io_Branch = _T_203 ? 1'h0 : _T_466; // @[control.py:97:Tile.fir@697.4]
  assign io_Branch_Src = _T_203 ? 1'h0 : _T_504; // @[control.py:98:Tile.fir@698.4]
  assign io_Mem_Read = _T_203 ? 1'h0 : _T_542; // @[control.py:102:Tile.fir@700.4]
  assign io_Mem_Write = _T_203 ? 1'h0 : _T_580; // @[control.py:103:Tile.fir@701.4]
  assign io_Data_Size = _T_203 ? 2'h0 : _T_618; // @[control.py:104:Tile.fir@702.4]
  assign io_Load_Type = _T_203 ? 1'h0 : _T_656; // @[control.py:105:Tile.fir@703.4]
  assign io_Mem_to_Reg = _T_203 ? 3'h0 : _T_694; // @[control.py:109:Tile.fir@705.4]
  assign io_Jump_Type = _T_203 ? 1'h0 : _T_732; // @[control.py:99:Tile.fir@699.4]
endmodule
module Tile( // @[tile.py:57:Tile.fir@708.2]
  input         clock, // @[rawmodule.py:100:Tile.fir@709.4]
  input         reset, // @[rawmodule.py:101:Tile.fir@710.4]
  input         io_PC_Write, // @[tile.py:18:Tile.fir@711.4]
  input  [31:0] io_pc_recover, // @[tile.py:18:Tile.fir@711.4]
  input  [31:0] io_new_addr, // @[tile.py:18:Tile.fir@711.4]
  input  [1:0]  io_PC_Sel, // @[tile.py:18:Tile.fir@711.4]
  input  [31:0] io_rd, // @[tile.py:18:Tile.fir@711.4]
  input  [31:0] io_wdata, // @[tile.py:18:Tile.fir@711.4]
  output        io_Reg_Write, // @[tile.py:18:Tile.fir@711.4]
  input         io_IF_ID_Write, // @[tile.py:18:Tile.fir@711.4]
  input         io_IF_ID_Flush, // @[tile.py:18:Tile.fir@711.4]
  output [2:0]  io_Imm_Sel, // @[tile.py:18:Tile.fir@711.4]
  output [31:0] io_id_pc, // @[tile.py:18:Tile.fir@711.4]
  output [31:0] io_id_pc_4, // @[tile.py:18:Tile.fir@711.4]
  output [31:0] io_id_inst, // @[tile.py:18:Tile.fir@711.4]
  output [31:0] io_rs1_out, // @[tile.py:18:Tile.fir@711.4]
  output [31:0] io_rs2_out, // @[tile.py:18:Tile.fir@711.4]
  output [31:0] io_imm, // @[tile.py:18:Tile.fir@711.4]
  output        io_ALU_Src, // @[tile.py:18:Tile.fir@711.4]
  output [4:0]  io_ALUOp, // @[tile.py:18:Tile.fir@711.4]
  output        io_Branch, // @[tile.py:18:Tile.fir@711.4]
  output        io_Branch_Src, // @[tile.py:18:Tile.fir@711.4]
  output        io_Mem_Read, // @[tile.py:18:Tile.fir@711.4]
  output        io_Mem_Write, // @[tile.py:18:Tile.fir@711.4]
  output [1:0]  io_Data_Size, // @[tile.py:18:Tile.fir@711.4]
  output        io_Load_Type, // @[tile.py:18:Tile.fir@711.4]
  output [2:0]  io_Mem_to_Reg, // @[tile.py:18:Tile.fir@711.4]
  output        io_Jump_Type // @[tile.py:18:Tile.fir@711.4]
);
  wire  pc_clock; // @[:Tile.fir@713.4]
  wire  pc_reset; // @[:Tile.fir@713.4]
  wire [31:0] pc_io_next_pc; // @[:Tile.fir@713.4]
  wire  pc_io_PC_Write; // @[:Tile.fir@713.4]
  wire [31:0] pc_io_pc_out; // @[:Tile.fir@713.4]
  wire  instcache_clock; // @[:Tile.fir@716.4]
  wire [31:0] instcache_io_addr; // @[:Tile.fir@716.4]
  wire [31:0] instcache_io_inst; // @[:Tile.fir@716.4]
  wire [31:0] datapath_io_if_io_pc_out; // @[:Tile.fir@719.4]
  wire [31:0] datapath_io_if_io_pc_recover; // @[:Tile.fir@719.4]
  wire [31:0] datapath_io_if_io_new_addr; // @[:Tile.fir@719.4]
  wire [31:0] datapath_io_if_io_next_pc; // @[:Tile.fir@719.4]
  wire [31:0] datapath_io_if_io_pc_4; // @[:Tile.fir@719.4]
  wire [1:0] datapath_io_if_io_PC_Sel; // @[:Tile.fir@719.4]
  wire  if_id_register_clock; // @[:Tile.fir@722.4]
  wire  if_id_register_reset; // @[:Tile.fir@722.4]
  wire [31:0] if_id_register_io_if_pc; // @[:Tile.fir@722.4]
  wire [31:0] if_id_register_io_if_pc_4; // @[:Tile.fir@722.4]
  wire [31:0] if_id_register_io_if_inst; // @[:Tile.fir@722.4]
  wire [31:0] if_id_register_io_id_pc; // @[:Tile.fir@722.4]
  wire [31:0] if_id_register_io_id_pc_4; // @[:Tile.fir@722.4]
  wire [4:0] if_id_register_io_id_rs1; // @[:Tile.fir@722.4]
  wire [4:0] if_id_register_io_id_rs2; // @[:Tile.fir@722.4]
  wire [31:0] if_id_register_io_id_inst; // @[:Tile.fir@722.4]
  wire  if_id_register_io_IF_ID_Write; // @[:Tile.fir@722.4]
  wire  if_id_register_io_IF_ID_Flush; // @[:Tile.fir@722.4]
  wire  regfile_clock; // @[:Tile.fir@725.4]
  wire [4:0] regfile_io_rs1; // @[:Tile.fir@725.4]
  wire [4:0] regfile_io_rs2; // @[:Tile.fir@725.4]
  wire [4:0] regfile_io_rd; // @[:Tile.fir@725.4]
  wire [31:0] regfile_io_wdata; // @[:Tile.fir@725.4]
  wire [31:0] regfile_io_rs1_out; // @[:Tile.fir@725.4]
  wire [31:0] regfile_io_rs2_out; // @[:Tile.fir@725.4]
  wire  regfile_io_Reg_Write; // @[:Tile.fir@725.4]
  wire [31:0] immgen_io_inst; // @[:Tile.fir@728.4]
  wire [31:0] immgen_io_imm; // @[:Tile.fir@728.4]
  wire [2:0] immgen_io_Imm_Sel; // @[:Tile.fir@728.4]
  wire [31:0] control_io_inst; // @[:Tile.fir@731.4]
  wire  control_io_Reg_Write; // @[:Tile.fir@731.4]
  wire [2:0] control_io_Imm_Sel; // @[:Tile.fir@731.4]
  wire  control_io_ALU_Src; // @[:Tile.fir@731.4]
  wire [4:0] control_io_ALUOp; // @[:Tile.fir@731.4]
  wire  control_io_Branch; // @[:Tile.fir@731.4]
  wire  control_io_Branch_Src; // @[:Tile.fir@731.4]
  wire  control_io_Mem_Read; // @[:Tile.fir@731.4]
  wire  control_io_Mem_Write; // @[:Tile.fir@731.4]
  wire [1:0] control_io_Data_Size; // @[:Tile.fir@731.4]
  wire  control_io_Load_Type; // @[:Tile.fir@731.4]
  wire [2:0] control_io_Mem_to_Reg; // @[:Tile.fir@731.4]
  wire  control_io_Jump_Type; // @[:Tile.fir@731.4]
  PC pc ( // @[:Tile.fir@713.4]
    .clock(pc_clock),
    .reset(pc_reset),
    .io_next_pc(pc_io_next_pc),
    .io_PC_Write(pc_io_PC_Write),
    .io_pc_out(pc_io_pc_out)
  );
  InstCache instcache ( // @[:Tile.fir@716.4]
    .clock(instcache_clock),
    .io_addr(instcache_io_addr),
    .io_inst(instcache_io_inst)
  );
  Datapath datapath ( // @[:Tile.fir@719.4]
    .io_if_io_pc_out(datapath_io_if_io_pc_out),
    .io_if_io_pc_recover(datapath_io_if_io_pc_recover),
    .io_if_io_new_addr(datapath_io_if_io_new_addr),
    .io_if_io_next_pc(datapath_io_if_io_next_pc),
    .io_if_io_pc_4(datapath_io_if_io_pc_4),
    .io_if_io_PC_Sel(datapath_io_if_io_PC_Sel)
  );
  IF_ID_Register if_id_register ( // @[:Tile.fir@722.4]
    .clock(if_id_register_clock),
    .reset(if_id_register_reset),
    .io_if_pc(if_id_register_io_if_pc),
    .io_if_pc_4(if_id_register_io_if_pc_4),
    .io_if_inst(if_id_register_io_if_inst),
    .io_id_pc(if_id_register_io_id_pc),
    .io_id_pc_4(if_id_register_io_id_pc_4),
    .io_id_rs1(if_id_register_io_id_rs1),
    .io_id_rs2(if_id_register_io_id_rs2),
    .io_id_inst(if_id_register_io_id_inst),
    .io_IF_ID_Write(if_id_register_io_IF_ID_Write),
    .io_IF_ID_Flush(if_id_register_io_IF_ID_Flush)
  );
  RegFile regfile ( // @[:Tile.fir@725.4]
    .clock(regfile_clock),
    .io_rs1(regfile_io_rs1),
    .io_rs2(regfile_io_rs2),
    .io_rd(regfile_io_rd),
    .io_wdata(regfile_io_wdata),
    .io_rs1_out(regfile_io_rs1_out),
    .io_rs2_out(regfile_io_rs2_out),
    .io_Reg_Write(regfile_io_Reg_Write)
  );
  ImmGen immgen ( // @[:Tile.fir@728.4]
    .io_inst(immgen_io_inst),
    .io_imm(immgen_io_imm),
    .io_Imm_Sel(immgen_io_Imm_Sel)
  );
  Control control ( // @[:Tile.fir@731.4]
    .io_inst(control_io_inst),
    .io_Reg_Write(control_io_Reg_Write),
    .io_Imm_Sel(control_io_Imm_Sel),
    .io_ALU_Src(control_io_ALU_Src),
    .io_ALUOp(control_io_ALUOp),
    .io_Branch(control_io_Branch),
    .io_Branch_Src(control_io_Branch_Src),
    .io_Mem_Read(control_io_Mem_Read),
    .io_Mem_Write(control_io_Mem_Write),
    .io_Data_Size(control_io_Data_Size),
    .io_Load_Type(control_io_Load_Type),
    .io_Mem_to_Reg(control_io_Mem_to_Reg),
    .io_Jump_Type(control_io_Jump_Type)
  );
  assign io_Reg_Write = control_io_Reg_Write; // @[tile.py:129:Tile.fir@760.4]
  assign io_Imm_Sel = control_io_Imm_Sel; // @[tile.py:130:Tile.fir@761.4]
  assign io_id_pc = if_id_register_io_id_pc; // @[tile.py:122:Tile.fir@754.4]
  assign io_id_pc_4 = if_id_register_io_id_pc_4; // @[tile.py:123:Tile.fir@755.4]
  assign io_id_inst = if_id_register_io_id_inst; // @[tile.py:124:Tile.fir@756.4]
  assign io_rs1_out = regfile_io_rs1_out; // @[tile.py:125:Tile.fir@757.4]
  assign io_rs2_out = regfile_io_rs2_out; // @[tile.py:126:Tile.fir@758.4]
  assign io_imm = immgen_io_imm; // @[tile.py:127:Tile.fir@759.4]
  assign io_ALU_Src = control_io_ALU_Src; // @[tile.py:131:Tile.fir@762.4]
  assign io_ALUOp = control_io_ALUOp; // @[tile.py:132:Tile.fir@763.4]
  assign io_Branch = control_io_Branch; // @[tile.py:133:Tile.fir@764.4]
  assign io_Branch_Src = control_io_Branch_Src; // @[tile.py:134:Tile.fir@765.4]
  assign io_Mem_Read = control_io_Mem_Read; // @[tile.py:135:Tile.fir@766.4]
  assign io_Mem_Write = control_io_Mem_Write; // @[tile.py:136:Tile.fir@767.4]
  assign io_Data_Size = control_io_Data_Size; // @[tile.py:137:Tile.fir@768.4]
  assign io_Load_Type = control_io_Load_Type; // @[tile.py:138:Tile.fir@769.4]
  assign io_Mem_to_Reg = control_io_Mem_to_Reg; // @[tile.py:139:Tile.fir@770.4]
  assign io_Jump_Type = control_io_Jump_Type; // @[tile.py:140:Tile.fir@771.4]
  assign pc_clock = clock; // @[rawmodule.py:110:Tile.fir@714.4]
  assign pc_reset = reset; // @[rawmodule.py:110:Tile.fir@715.4]
  assign pc_io_next_pc = datapath_io_if_io_next_pc; // @[tile.py:74:Tile.fir@734.4]
  assign pc_io_PC_Write = io_PC_Write; // @[tile.py:75:Tile.fir@735.4]
  assign instcache_clock = clock; // @[rawmodule.py:110:Tile.fir@717.4]
  assign instcache_io_addr = pc_io_pc_out; // @[tile.py:80:Tile.fir@736.4]
  assign datapath_io_if_io_pc_out = pc_io_pc_out; // @[tile.py:85:Tile.fir@737.4]
  assign datapath_io_if_io_pc_recover = io_pc_recover; // @[tile.py:86:Tile.fir@738.4]
  assign datapath_io_if_io_new_addr = io_new_addr; // @[tile.py:87:Tile.fir@739.4]
  assign datapath_io_if_io_PC_Sel = io_PC_Sel; // @[tile.py:88:Tile.fir@740.4]
  assign if_id_register_clock = clock; // @[rawmodule.py:110:Tile.fir@723.4]
  assign if_id_register_reset = reset; // @[rawmodule.py:110:Tile.fir@724.4]
  assign if_id_register_io_if_pc = pc_io_pc_out; // @[tile.py:93:Tile.fir@741.4]
  assign if_id_register_io_if_pc_4 = datapath_io_if_io_pc_4; // @[tile.py:94:Tile.fir@742.4]
  assign if_id_register_io_if_inst = instcache_io_inst; // @[tile.py:95:Tile.fir@743.4]
  assign if_id_register_io_IF_ID_Write = io_IF_ID_Write; // @[tile.py:97:Tile.fir@745.4]
  assign if_id_register_io_IF_ID_Flush = io_IF_ID_Flush; // @[tile.py:96:Tile.fir@744.4]
  assign regfile_clock = clock; // @[rawmodule.py:110:Tile.fir@726.4]
  assign regfile_io_rs1 = if_id_register_io_id_rs1; // @[tile.py:102:Tile.fir@746.4]
  assign regfile_io_rs2 = if_id_register_io_id_rs2; // @[tile.py:103:Tile.fir@747.4]
  assign regfile_io_rd = io_rd[4:0]; // @[tile.py:104:Tile.fir@748.4]
  assign regfile_io_wdata = io_wdata; // @[tile.py:105:Tile.fir@749.4]
  assign regfile_io_Reg_Write = control_io_Reg_Write; // @[tile.py:106:Tile.fir@750.4]
  assign immgen_io_inst = if_id_register_io_id_inst; // @[tile.py:111:Tile.fir@751.4]
  assign immgen_io_Imm_Sel = control_io_Imm_Sel; // @[tile.py:112:Tile.fir@752.4]
  assign control_io_inst = if_id_register_io_id_inst; // @[tile.py:117:Tile.fir@753.4]
endmodule
